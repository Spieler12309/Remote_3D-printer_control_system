module delay(
input 	wire 				clk,
input		wire	[31:0]	delay,

output	wire				done



endmodule
