module find_max_timing(	
	input		wire				clk,
	input		wire				reset,
	input		wire				start,
	input		wire	[31:0]	params_a [0:4],
	input		wire	[31:0]	params_b [0:4],
	input		wire	[31:0]	params_z [0:4],
	input		wire	[31:0]	params_e [0:4],
	
	input		wire	[63:0]	timing_a	[0:3],
	input		wire	[63:0]	timing_b	[0:3],
	input		wire	[63:0]	timing_z	[0:3],
	input		wire	[63:0]	timing_e	[0:3],


	output	wire	[63:0]	max_timing 	[0:3],
	output	reg				finish	
	);

endmodule
