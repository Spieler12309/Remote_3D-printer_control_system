// soc_system.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module soc_system (
		input  wire        clk_clk,                                             //                                          clk.clk
		output wire [11:0] command_dt_external_connection_export,               //               command_dt_external_connection.export
		output wire [31:0] command_e0_external_connection_export,               //               command_e0_external_connection.export
		output wire [31:0] command_e1_external_connection_export,               //               command_e1_external_connection.export
		output wire [31:0] command_f_e0_external_connection_export,             //             command_f_e0_external_connection.export
		output wire [31:0] command_f_e1_external_connection_export,             //             command_f_e1_external_connection.export
		output wire [31:0] command_f_x_external_connection_export,              //              command_f_x_external_connection.export
		output wire [31:0] command_f_y_external_connection_export,              //              command_f_y_external_connection.export
		output wire [31:0] command_f_z_external_connection_export,              //              command_f_z_external_connection.export
		output wire [11:0] command_t_external_connection_export,                //                command_t_external_connection.export
		output wire [31:0] command_type_external_connection_export,             //             command_type_external_connection.export
		output wire [31:0] command_x_external_connection_export,                //                command_x_external_connection.export
		output wire [31:0] command_y_external_connection_export,                //                command_y_external_connection.export
		output wire [31:0] command_z_external_connection_export,                //                command_z_external_connection.export
		input  wire [31:0] flags_in_external_connection_export,                 //                 flags_in_external_connection.export
		output wire [31:0] flags_out_external_connection_export,                //                flags_out_external_connection.export
		input  wire        hps_0_f2h_cold_reset_req_reset_n,                    //                     hps_0_f2h_cold_reset_req.reset_n
		input  wire        hps_0_f2h_debug_reset_req_reset_n,                   //                    hps_0_f2h_debug_reset_req.reset_n
		input  wire [27:0] hps_0_f2h_stm_hw_events_stm_hwevents,                //                      hps_0_f2h_stm_hw_events.stm_hwevents
		input  wire        hps_0_f2h_warm_reset_req_reset_n,                    //                     hps_0_f2h_warm_reset_req.reset_n
		output wire        hps_0_h2f_reset_reset_n,                             //                              hps_0_h2f_reset.reset_n
		output wire        hps_0_hps_io_hps_io_emac1_inst_TX_CLK,               //                                 hps_0_hps_io.hps_io_emac1_inst_TX_CLK
		output wire        hps_0_hps_io_hps_io_emac1_inst_TXD0,                 //                                             .hps_io_emac1_inst_TXD0
		output wire        hps_0_hps_io_hps_io_emac1_inst_TXD1,                 //                                             .hps_io_emac1_inst_TXD1
		output wire        hps_0_hps_io_hps_io_emac1_inst_TXD2,                 //                                             .hps_io_emac1_inst_TXD2
		output wire        hps_0_hps_io_hps_io_emac1_inst_TXD3,                 //                                             .hps_io_emac1_inst_TXD3
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RXD0,                 //                                             .hps_io_emac1_inst_RXD0
		inout  wire        hps_0_hps_io_hps_io_emac1_inst_MDIO,                 //                                             .hps_io_emac1_inst_MDIO
		output wire        hps_0_hps_io_hps_io_emac1_inst_MDC,                  //                                             .hps_io_emac1_inst_MDC
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RX_CTL,               //                                             .hps_io_emac1_inst_RX_CTL
		output wire        hps_0_hps_io_hps_io_emac1_inst_TX_CTL,               //                                             .hps_io_emac1_inst_TX_CTL
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RX_CLK,               //                                             .hps_io_emac1_inst_RX_CLK
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RXD1,                 //                                             .hps_io_emac1_inst_RXD1
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RXD2,                 //                                             .hps_io_emac1_inst_RXD2
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RXD3,                 //                                             .hps_io_emac1_inst_RXD3
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_CMD,                   //                                             .hps_io_sdio_inst_CMD
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_D0,                    //                                             .hps_io_sdio_inst_D0
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_D1,                    //                                             .hps_io_sdio_inst_D1
		output wire        hps_0_hps_io_hps_io_sdio_inst_CLK,                   //                                             .hps_io_sdio_inst_CLK
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_D2,                    //                                             .hps_io_sdio_inst_D2
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_D3,                    //                                             .hps_io_sdio_inst_D3
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D0,                    //                                             .hps_io_usb1_inst_D0
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D1,                    //                                             .hps_io_usb1_inst_D1
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D2,                    //                                             .hps_io_usb1_inst_D2
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D3,                    //                                             .hps_io_usb1_inst_D3
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D4,                    //                                             .hps_io_usb1_inst_D4
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D5,                    //                                             .hps_io_usb1_inst_D5
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D6,                    //                                             .hps_io_usb1_inst_D6
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D7,                    //                                             .hps_io_usb1_inst_D7
		input  wire        hps_0_hps_io_hps_io_usb1_inst_CLK,                   //                                             .hps_io_usb1_inst_CLK
		output wire        hps_0_hps_io_hps_io_usb1_inst_STP,                   //                                             .hps_io_usb1_inst_STP
		input  wire        hps_0_hps_io_hps_io_usb1_inst_DIR,                   //                                             .hps_io_usb1_inst_DIR
		input  wire        hps_0_hps_io_hps_io_usb1_inst_NXT,                   //                                             .hps_io_usb1_inst_NXT
		output wire        hps_0_hps_io_hps_io_spim1_inst_CLK,                  //                                             .hps_io_spim1_inst_CLK
		output wire        hps_0_hps_io_hps_io_spim1_inst_MOSI,                 //                                             .hps_io_spim1_inst_MOSI
		input  wire        hps_0_hps_io_hps_io_spim1_inst_MISO,                 //                                             .hps_io_spim1_inst_MISO
		output wire        hps_0_hps_io_hps_io_spim1_inst_SS0,                  //                                             .hps_io_spim1_inst_SS0
		input  wire        hps_0_hps_io_hps_io_uart0_inst_RX,                   //                                             .hps_io_uart0_inst_RX
		output wire        hps_0_hps_io_hps_io_uart0_inst_TX,                   //                                             .hps_io_uart0_inst_TX
		inout  wire        hps_0_hps_io_hps_io_i2c0_inst_SDA,                   //                                             .hps_io_i2c0_inst_SDA
		inout  wire        hps_0_hps_io_hps_io_i2c0_inst_SCL,                   //                                             .hps_io_i2c0_inst_SCL
		inout  wire        hps_0_hps_io_hps_io_i2c1_inst_SDA,                   //                                             .hps_io_i2c1_inst_SDA
		inout  wire        hps_0_hps_io_hps_io_i2c1_inst_SCL,                   //                                             .hps_io_i2c1_inst_SCL
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO09,                //                                             .hps_io_gpio_inst_GPIO09
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO35,                //                                             .hps_io_gpio_inst_GPIO35
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO40,                //                                             .hps_io_gpio_inst_GPIO40
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO53,                //                                             .hps_io_gpio_inst_GPIO53
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO54,                //                                             .hps_io_gpio_inst_GPIO54
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO61,                //                                             .hps_io_gpio_inst_GPIO61
		input  wire        hps_0_uart1_cts,                                     //                                  hps_0_uart1.cts
		input  wire        hps_0_uart1_dsr,                                     //                                             .dsr
		input  wire        hps_0_uart1_dcd,                                     //                                             .dcd
		input  wire        hps_0_uart1_ri,                                      //                                             .ri
		output wire        hps_0_uart1_dtr,                                     //                                             .dtr
		output wire        hps_0_uart1_rts,                                     //                                             .rts
		output wire        hps_0_uart1_out1_n,                                  //                                             .out1_n
		output wire        hps_0_uart1_out2_n,                                  //                                             .out2_n
		input  wire        hps_0_uart1_rxd,                                     //                                             .rxd
		output wire        hps_0_uart1_txd,                                     //                                             .txd
		input  wire [31:0] max_params_0_external_connection_export,             //             max_params_0_external_connection.export
		input  wire [31:0] max_params_1_external_connection_export,             //             max_params_1_external_connection.export
		input  wire [31:0] max_params_2_external_connection_export,             //             max_params_2_external_connection.export
		input  wire [31:0] max_params_3_external_connection_export,             //             max_params_3_external_connection.export
		input  wire [31:0] max_params_4_external_connection_export,             //             max_params_4_external_connection.export
		input  wire [31:0] max_timing_0_external_connection_export,             //             max_timing_0_external_connection.export
		input  wire [31:0] max_timing_1_external_connection_export,             //             max_timing_1_external_connection.export
		input  wire [31:0] max_timing_2_external_connection_export,             //             max_timing_2_external_connection.export
		input  wire [31:0] max_timing_3_external_connection_export,             //             max_timing_3_external_connection.export
		output wire [14:0] memory_mem_a,                                        //                                       memory.mem_a
		output wire [2:0]  memory_mem_ba,                                       //                                             .mem_ba
		output wire        memory_mem_ck,                                       //                                             .mem_ck
		output wire        memory_mem_ck_n,                                     //                                             .mem_ck_n
		output wire        memory_mem_cke,                                      //                                             .mem_cke
		output wire        memory_mem_cs_n,                                     //                                             .mem_cs_n
		output wire        memory_mem_ras_n,                                    //                                             .mem_ras_n
		output wire        memory_mem_cas_n,                                    //                                             .mem_cas_n
		output wire        memory_mem_we_n,                                     //                                             .mem_we_n
		output wire        memory_mem_reset_n,                                  //                                             .mem_reset_n
		inout  wire [31:0] memory_mem_dq,                                       //                                             .mem_dq
		inout  wire [3:0]  memory_mem_dqs,                                      //                                             .mem_dqs
		inout  wire [3:0]  memory_mem_dqs_n,                                    //                                             .mem_dqs_n
		output wire        memory_mem_odt,                                      //                                             .mem_odt
		output wire [3:0]  memory_mem_dm,                                       //                                             .mem_dm
		input  wire        memory_oct_rzqin,                                    //                                             .oct_rzqin
		input  wire [31:0] new_rparams_e0_0_external_connection_export,         //         new_rparams_e0_0_external_connection.export
		input  wire [31:0] new_rparams_e0_1_external_connection_export,         //         new_rparams_e0_1_external_connection.export
		input  wire [31:0] new_rparams_e0_2_external_connection_export,         //         new_rparams_e0_2_external_connection.export
		input  wire [31:0] new_rparams_e0_3_external_connection_export,         //         new_rparams_e0_3_external_connection.export
		input  wire [31:0] new_rparams_e0_4_external_connection_export,         //         new_rparams_e0_4_external_connection.export
		input  wire [31:0] new_rparams_e1_0_external_connection_export,         //         new_rparams_e1_0_external_connection.export
		input  wire [31:0] new_rparams_e1_1_external_connection_export,         //         new_rparams_e1_1_external_connection.export
		input  wire [31:0] new_rparams_e1_2_external_connection_export,         //         new_rparams_e1_2_external_connection.export
		input  wire [31:0] new_rparams_e1_3_external_connection_export,         //         new_rparams_e1_3_external_connection.export
		input  wire [31:0] new_rparams_e1_4_external_connection_export,         //         new_rparams_e1_4_external_connection.export
		input  wire [31:0] new_rparams_x_0_external_connection_export,          //          new_rparams_x_0_external_connection.export
		input  wire [31:0] new_rparams_x_1_external_connection_export,          //          new_rparams_x_1_external_connection.export
		input  wire [31:0] new_rparams_x_2_external_connection_export,          //          new_rparams_x_2_external_connection.export
		input  wire [31:0] new_rparams_x_3_external_connection_export,          //          new_rparams_x_3_external_connection.export
		input  wire [31:0] new_rparams_x_4_external_connection_export,          //          new_rparams_x_4_external_connection.export
		input  wire [31:0] new_rparams_y_0_external_connection_export,          //          new_rparams_y_0_external_connection.export
		input  wire [31:0] new_rparams_y_1_external_connection_export,          //          new_rparams_y_1_external_connection.export
		input  wire [31:0] new_rparams_y_2_external_connection_export,          //          new_rparams_y_2_external_connection.export
		input  wire [31:0] new_rparams_y_3_external_connection_export,          //          new_rparams_y_3_external_connection.export
		input  wire [31:0] new_rparams_y_4_external_connection_export,          //          new_rparams_y_4_external_connection.export
		input  wire [31:0] new_rparams_z_0_external_connection_export,          //          new_rparams_z_0_external_connection.export
		input  wire [31:0] new_rparams_z_1_external_connection_export,          //          new_rparams_z_1_external_connection.export
		input  wire [31:0] new_rparams_z_2_external_connection_export,          //          new_rparams_z_2_external_connection.export
		input  wire [31:0] new_rparams_z_3_external_connection_export,          //          new_rparams_z_3_external_connection.export
		input  wire [31:0] new_rparams_z_4_external_connection_export,          //          new_rparams_z_4_external_connection.export
		input  wire [31:0] params_e0_0_external_connection_export,              //              params_e0_0_external_connection.export
		input  wire [31:0] params_e0_1_external_connection_export,              //              params_e0_1_external_connection.export
		input  wire [31:0] params_e0_2_external_connection_export,              //              params_e0_2_external_connection.export
		input  wire [31:0] params_e0_3_external_connection_export,              //              params_e0_3_external_connection.export
		input  wire [31:0] params_e0_4_external_connection_export,              //              params_e0_4_external_connection.export
		input  wire [31:0] params_e1_0_external_connection_export,              //              params_e1_0_external_connection.export
		input  wire [31:0] params_e1_1_external_connection_export,              //              params_e1_1_external_connection.export
		input  wire [31:0] params_e1_2_external_connection_export,              //              params_e1_2_external_connection.export
		input  wire [31:0] params_e1_3_external_connection_export,              //              params_e1_3_external_connection.export
		input  wire [31:0] params_e1_4_external_connection_export,              //              params_e1_4_external_connection.export
		input  wire [31:0] params_x_0_external_connection_export,               //               params_x_0_external_connection.export
		input  wire [31:0] params_x_1_external_connection_export,               //               params_x_1_external_connection.export
		input  wire [31:0] params_x_2_external_connection_export,               //               params_x_2_external_connection.export
		input  wire [31:0] params_x_3_external_connection_export,               //               params_x_3_external_connection.export
		input  wire [31:0] params_x_4_external_connection_export,               //               params_x_4_external_connection.export
		input  wire [31:0] params_y_0_external_connection_export,               //               params_y_0_external_connection.export
		input  wire [31:0] params_y_1_external_connection_export,               //               params_y_1_external_connection.export
		input  wire [31:0] params_y_2_external_connection_export,               //               params_y_2_external_connection.export
		input  wire [31:0] params_y_3_external_connection_export,               //               params_y_3_external_connection.export
		input  wire [31:0] params_y_4_external_connection_export,               //               params_y_4_external_connection.export
		input  wire [31:0] params_z_0_external_connection_export,               //               params_z_0_external_connection.export
		input  wire [31:0] params_z_1_external_connection_export,               //               params_z_1_external_connection.export
		input  wire [31:0] params_z_2_external_connection_export,               //               params_z_2_external_connection.export
		input  wire [31:0] params_z_3_external_connection_export,               //               params_z_3_external_connection.export
		input  wire [31:0] params_z_4_external_connection_export,               //               params_z_4_external_connection.export
		output wire        pll_sys_outclk100mhz_clk,                            //                         pll_sys_outclk100mhz.clk
		output wire        pll_sys_outclk10mhz_clk,                             //                          pll_sys_outclk10mhz.clk
		output wire        pll_sys_outclk1mhz_clk,                              //                           pll_sys_outclk1mhz.clk
		output wire        pll_sys_outclk5mhz_clk,                              //                           pll_sys_outclk5mhz.clk
		input  wire [11:0] position_e0_external_connection_export,              //              position_e0_external_connection.export
		input  wire [11:0] position_e1_external_connection_export,              //              position_e1_external_connection.export
		input  wire [11:0] position_x_external_connection_export,               //               position_x_external_connection.export
		input  wire [11:0] position_y_external_connection_export,               //               position_y_external_connection.export
		input  wire [11:0] position_z_external_connection_export,               //               position_z_external_connection.export
		input  wire        reset_reset_n,                                       //                                        reset.reset_n
		output wire [31:0] settings_acceleration_e0_external_connection_export, // settings_acceleration_e0_external_connection.export
		output wire [31:0] settings_acceleration_e1_external_connection_export, // settings_acceleration_e1_external_connection.export
		output wire [31:0] settings_acceleration_x_external_connection_export,  //  settings_acceleration_x_external_connection.export
		output wire [31:0] settings_acceleration_y_external_connection_export,  //  settings_acceleration_y_external_connection.export
		output wire [31:0] settings_acceleration_z_external_connection_export,  //  settings_acceleration_z_external_connection.export
		output wire [31:0] settings_jerk_e0_external_connection_export,         //         settings_jerk_e0_external_connection.export
		output wire [31:0] settings_jerk_e1_external_connection_export,         //         settings_jerk_e1_external_connection.export
		output wire [31:0] settings_jerk_x_external_connection_export,          //          settings_jerk_x_external_connection.export
		output wire [31:0] settings_jerk_y_external_connection_export,          //          settings_jerk_y_external_connection.export
		output wire [31:0] settings_jerk_z_external_connection_export,          //          settings_jerk_z_external_connection.export
		output wire [31:0] settings_max_speed_e0_external_connection_export,    //    settings_max_speed_e0_external_connection.export
		output wire [31:0] settings_max_speed_e1_external_connection_export,    //    settings_max_speed_e1_external_connection.export
		output wire [31:0] settings_max_speed_x_external_connection_export,     //     settings_max_speed_x_external_connection.export
		output wire [31:0] settings_max_speed_y_external_connection_export,     //     settings_max_speed_y_external_connection.export
		output wire [31:0] settings_max_speed_z_external_connection_export,     //     settings_max_speed_z_external_connection.export
		output wire [11:0] settings_max_temp_bed_external_connection_export,    //    settings_max_temp_bed_external_connection.export
		output wire [11:0] settings_max_temp_e0_external_connection_export,     //     settings_max_temp_e0_external_connection.export
		output wire [11:0] settings_max_temp_e1_external_connection_export,     //     settings_max_temp_e1_external_connection.export
		input  wire [31:0] step_e0_now_external_connection_export,              //              step_e0_now_external_connection.export
		input  wire [31:0] step_e1_now_external_connection_export,              //              step_e1_now_external_connection.export
		input  wire [31:0] step_x_now_external_connection_export,               //               step_x_now_external_connection.export
		input  wire [31:0] step_y_now_external_connection_export,               //               step_y_now_external_connection.export
		input  wire [31:0] step_z_now_external_connection_export,               //               step_z_now_external_connection.export
		input  wire [11:0] temp_0_external_connection_export,                   //                   temp_0_external_connection.export
		input  wire [11:0] temp_1_external_connection_export,                   //                   temp_1_external_connection.export
		input  wire [11:0] temp_2_external_connection_export,                   //                   temp_2_external_connection.export
		input  wire [31:0] timing_e0_0_external_connection_export,              //              timing_e0_0_external_connection.export
		input  wire [31:0] timing_e0_1_external_connection_export,              //              timing_e0_1_external_connection.export
		input  wire [31:0] timing_e0_2_external_connection_export,              //              timing_e0_2_external_connection.export
		input  wire [31:0] timing_e0_3_external_connection_export,              //              timing_e0_3_external_connection.export
		input  wire [31:0] timing_e1_0_external_connection_export,              //              timing_e1_0_external_connection.export
		input  wire [31:0] timing_e1_1_external_connection_export,              //              timing_e1_1_external_connection.export
		input  wire [31:0] timing_e1_2_external_connection_export,              //              timing_e1_2_external_connection.export
		input  wire [31:0] timing_e1_3_external_connection_export,              //              timing_e1_3_external_connection.export
		input  wire [31:0] timing_x_0_external_connection_export,               //               timing_x_0_external_connection.export
		input  wire [31:0] timing_x_1_external_connection_export,               //               timing_x_1_external_connection.export
		input  wire [31:0] timing_x_2_external_connection_export,               //               timing_x_2_external_connection.export
		input  wire [31:0] timing_x_3_external_connection_export,               //               timing_x_3_external_connection.export
		input  wire [31:0] timing_y_0_external_connection_export,               //               timing_y_0_external_connection.export
		input  wire [31:0] timing_y_1_external_connection_export,               //               timing_y_1_external_connection.export
		input  wire [31:0] timing_y_2_external_connection_export,               //               timing_y_2_external_connection.export
		input  wire [31:0] timing_y_3_external_connection_export,               //               timing_y_3_external_connection.export
		input  wire [31:0] timing_z_0_external_connection_export,               //               timing_z_0_external_connection.export
		input  wire [31:0] timing_z_1_external_connection_export,               //               timing_z_1_external_connection.export
		input  wire [31:0] timing_z_2_external_connection_export,               //               timing_z_2_external_connection.export
		input  wire [31:0] timing_z_3_external_connection_export                //               timing_z_3_external_connection.export
	);

	wire    [1:0] hps_0_h2f_lw_axi_master_awburst;                           // hps_0:h2f_lw_AWBURST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awburst
	wire    [3:0] hps_0_h2f_lw_axi_master_arlen;                             // hps_0:h2f_lw_ARLEN -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arlen
	wire    [3:0] hps_0_h2f_lw_axi_master_wstrb;                             // hps_0:h2f_lw_WSTRB -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wstrb
	wire          hps_0_h2f_lw_axi_master_wready;                            // mm_interconnect_0:hps_0_h2f_lw_axi_master_wready -> hps_0:h2f_lw_WREADY
	wire   [11:0] hps_0_h2f_lw_axi_master_rid;                               // mm_interconnect_0:hps_0_h2f_lw_axi_master_rid -> hps_0:h2f_lw_RID
	wire          hps_0_h2f_lw_axi_master_rready;                            // hps_0:h2f_lw_RREADY -> mm_interconnect_0:hps_0_h2f_lw_axi_master_rready
	wire    [3:0] hps_0_h2f_lw_axi_master_awlen;                             // hps_0:h2f_lw_AWLEN -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awlen
	wire   [11:0] hps_0_h2f_lw_axi_master_wid;                               // hps_0:h2f_lw_WID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wid
	wire    [3:0] hps_0_h2f_lw_axi_master_arcache;                           // hps_0:h2f_lw_ARCACHE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arcache
	wire          hps_0_h2f_lw_axi_master_wvalid;                            // hps_0:h2f_lw_WVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wvalid
	wire   [20:0] hps_0_h2f_lw_axi_master_araddr;                            // hps_0:h2f_lw_ARADDR -> mm_interconnect_0:hps_0_h2f_lw_axi_master_araddr
	wire    [2:0] hps_0_h2f_lw_axi_master_arprot;                            // hps_0:h2f_lw_ARPROT -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arprot
	wire    [2:0] hps_0_h2f_lw_axi_master_awprot;                            // hps_0:h2f_lw_AWPROT -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awprot
	wire   [31:0] hps_0_h2f_lw_axi_master_wdata;                             // hps_0:h2f_lw_WDATA -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wdata
	wire          hps_0_h2f_lw_axi_master_arvalid;                           // hps_0:h2f_lw_ARVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arvalid
	wire    [3:0] hps_0_h2f_lw_axi_master_awcache;                           // hps_0:h2f_lw_AWCACHE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awcache
	wire   [11:0] hps_0_h2f_lw_axi_master_arid;                              // hps_0:h2f_lw_ARID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arid
	wire    [1:0] hps_0_h2f_lw_axi_master_arlock;                            // hps_0:h2f_lw_ARLOCK -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arlock
	wire    [1:0] hps_0_h2f_lw_axi_master_awlock;                            // hps_0:h2f_lw_AWLOCK -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awlock
	wire   [20:0] hps_0_h2f_lw_axi_master_awaddr;                            // hps_0:h2f_lw_AWADDR -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awaddr
	wire    [1:0] hps_0_h2f_lw_axi_master_bresp;                             // mm_interconnect_0:hps_0_h2f_lw_axi_master_bresp -> hps_0:h2f_lw_BRESP
	wire          hps_0_h2f_lw_axi_master_arready;                           // mm_interconnect_0:hps_0_h2f_lw_axi_master_arready -> hps_0:h2f_lw_ARREADY
	wire   [31:0] hps_0_h2f_lw_axi_master_rdata;                             // mm_interconnect_0:hps_0_h2f_lw_axi_master_rdata -> hps_0:h2f_lw_RDATA
	wire          hps_0_h2f_lw_axi_master_awready;                           // mm_interconnect_0:hps_0_h2f_lw_axi_master_awready -> hps_0:h2f_lw_AWREADY
	wire    [1:0] hps_0_h2f_lw_axi_master_arburst;                           // hps_0:h2f_lw_ARBURST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arburst
	wire    [2:0] hps_0_h2f_lw_axi_master_arsize;                            // hps_0:h2f_lw_ARSIZE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arsize
	wire          hps_0_h2f_lw_axi_master_bready;                            // hps_0:h2f_lw_BREADY -> mm_interconnect_0:hps_0_h2f_lw_axi_master_bready
	wire          hps_0_h2f_lw_axi_master_rlast;                             // mm_interconnect_0:hps_0_h2f_lw_axi_master_rlast -> hps_0:h2f_lw_RLAST
	wire          hps_0_h2f_lw_axi_master_wlast;                             // hps_0:h2f_lw_WLAST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wlast
	wire    [1:0] hps_0_h2f_lw_axi_master_rresp;                             // mm_interconnect_0:hps_0_h2f_lw_axi_master_rresp -> hps_0:h2f_lw_RRESP
	wire   [11:0] hps_0_h2f_lw_axi_master_awid;                              // hps_0:h2f_lw_AWID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awid
	wire   [11:0] hps_0_h2f_lw_axi_master_bid;                               // mm_interconnect_0:hps_0_h2f_lw_axi_master_bid -> hps_0:h2f_lw_BID
	wire          hps_0_h2f_lw_axi_master_bvalid;                            // mm_interconnect_0:hps_0_h2f_lw_axi_master_bvalid -> hps_0:h2f_lw_BVALID
	wire    [2:0] hps_0_h2f_lw_axi_master_awsize;                            // hps_0:h2f_lw_AWSIZE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awsize
	wire          hps_0_h2f_lw_axi_master_awvalid;                           // hps_0:h2f_lw_AWVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awvalid
	wire          hps_0_h2f_lw_axi_master_rvalid;                            // mm_interconnect_0:hps_0_h2f_lw_axi_master_rvalid -> hps_0:h2f_lw_RVALID
	wire   [31:0] mm_interconnect_0_mm_bridge_0_s0_readdata;                 // mm_bridge_0:s0_readdata -> mm_interconnect_0:mm_bridge_0_s0_readdata
	wire          mm_interconnect_0_mm_bridge_0_s0_waitrequest;              // mm_bridge_0:s0_waitrequest -> mm_interconnect_0:mm_bridge_0_s0_waitrequest
	wire          mm_interconnect_0_mm_bridge_0_s0_debugaccess;              // mm_interconnect_0:mm_bridge_0_s0_debugaccess -> mm_bridge_0:s0_debugaccess
	wire   [17:0] mm_interconnect_0_mm_bridge_0_s0_address;                  // mm_interconnect_0:mm_bridge_0_s0_address -> mm_bridge_0:s0_address
	wire          mm_interconnect_0_mm_bridge_0_s0_read;                     // mm_interconnect_0:mm_bridge_0_s0_read -> mm_bridge_0:s0_read
	wire    [3:0] mm_interconnect_0_mm_bridge_0_s0_byteenable;               // mm_interconnect_0:mm_bridge_0_s0_byteenable -> mm_bridge_0:s0_byteenable
	wire          mm_interconnect_0_mm_bridge_0_s0_readdatavalid;            // mm_bridge_0:s0_readdatavalid -> mm_interconnect_0:mm_bridge_0_s0_readdatavalid
	wire          mm_interconnect_0_mm_bridge_0_s0_write;                    // mm_interconnect_0:mm_bridge_0_s0_write -> mm_bridge_0:s0_write
	wire   [31:0] mm_interconnect_0_mm_bridge_0_s0_writedata;                // mm_interconnect_0:mm_bridge_0_s0_writedata -> mm_bridge_0:s0_writedata
	wire    [0:0] mm_interconnect_0_mm_bridge_0_s0_burstcount;               // mm_interconnect_0:mm_bridge_0_s0_burstcount -> mm_bridge_0:s0_burstcount
	wire          mm_bridge_0_m0_waitrequest;                                // mm_interconnect_1:mm_bridge_0_m0_waitrequest -> mm_bridge_0:m0_waitrequest
	wire   [31:0] mm_bridge_0_m0_readdata;                                   // mm_interconnect_1:mm_bridge_0_m0_readdata -> mm_bridge_0:m0_readdata
	wire          mm_bridge_0_m0_debugaccess;                                // mm_bridge_0:m0_debugaccess -> mm_interconnect_1:mm_bridge_0_m0_debugaccess
	wire   [17:0] mm_bridge_0_m0_address;                                    // mm_bridge_0:m0_address -> mm_interconnect_1:mm_bridge_0_m0_address
	wire          mm_bridge_0_m0_read;                                       // mm_bridge_0:m0_read -> mm_interconnect_1:mm_bridge_0_m0_read
	wire    [3:0] mm_bridge_0_m0_byteenable;                                 // mm_bridge_0:m0_byteenable -> mm_interconnect_1:mm_bridge_0_m0_byteenable
	wire          mm_bridge_0_m0_readdatavalid;                              // mm_interconnect_1:mm_bridge_0_m0_readdatavalid -> mm_bridge_0:m0_readdatavalid
	wire   [31:0] mm_bridge_0_m0_writedata;                                  // mm_bridge_0:m0_writedata -> mm_interconnect_1:mm_bridge_0_m0_writedata
	wire          mm_bridge_0_m0_write;                                      // mm_bridge_0:m0_write -> mm_interconnect_1:mm_bridge_0_m0_write
	wire    [0:0] mm_bridge_0_m0_burstcount;                                 // mm_bridge_0:m0_burstcount -> mm_interconnect_1:mm_bridge_0_m0_burstcount
	wire   [31:0] fpga_only_master_master_readdata;                          // mm_interconnect_1:fpga_only_master_master_readdata -> fpga_only_master:master_readdata
	wire          fpga_only_master_master_waitrequest;                       // mm_interconnect_1:fpga_only_master_master_waitrequest -> fpga_only_master:master_waitrequest
	wire   [31:0] fpga_only_master_master_address;                           // fpga_only_master:master_address -> mm_interconnect_1:fpga_only_master_master_address
	wire          fpga_only_master_master_read;                              // fpga_only_master:master_read -> mm_interconnect_1:fpga_only_master_master_read
	wire    [3:0] fpga_only_master_master_byteenable;                        // fpga_only_master:master_byteenable -> mm_interconnect_1:fpga_only_master_master_byteenable
	wire          fpga_only_master_master_readdatavalid;                     // mm_interconnect_1:fpga_only_master_master_readdatavalid -> fpga_only_master:master_readdatavalid
	wire          fpga_only_master_master_write;                             // fpga_only_master:master_write -> mm_interconnect_1:fpga_only_master_master_write
	wire   [31:0] fpga_only_master_master_writedata;                         // fpga_only_master:master_writedata -> mm_interconnect_1:fpga_only_master_master_writedata
	wire          mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect;  // mm_interconnect_1:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire   [31:0] mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata;    // jtag_uart:av_readdata -> mm_interconnect_1:jtag_uart_avalon_jtag_slave_readdata
	wire          mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest; // jtag_uart:av_waitrequest -> mm_interconnect_1:jtag_uart_avalon_jtag_slave_waitrequest
	wire    [0:0] mm_interconnect_1_jtag_uart_avalon_jtag_slave_address;     // mm_interconnect_1:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire          mm_interconnect_1_jtag_uart_avalon_jtag_slave_read;        // mm_interconnect_1:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire          mm_interconnect_1_jtag_uart_avalon_jtag_slave_write;       // mm_interconnect_1:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire   [31:0] mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata;   // mm_interconnect_1:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire   [31:0] mm_interconnect_1_ilc_avalon_slave_readdata;               // ILC:avmm_rddata -> mm_interconnect_1:ILC_avalon_slave_readdata
	wire    [5:0] mm_interconnect_1_ilc_avalon_slave_address;                // mm_interconnect_1:ILC_avalon_slave_address -> ILC:avmm_addr
	wire          mm_interconnect_1_ilc_avalon_slave_read;                   // mm_interconnect_1:ILC_avalon_slave_read -> ILC:avmm_read
	wire          mm_interconnect_1_ilc_avalon_slave_write;                  // mm_interconnect_1:ILC_avalon_slave_write -> ILC:avmm_write
	wire   [31:0] mm_interconnect_1_ilc_avalon_slave_writedata;              // mm_interconnect_1:ILC_avalon_slave_writedata -> ILC:avmm_wrdata
	wire   [31:0] mm_interconnect_1_sysid_qsys_control_slave_readdata;       // sysid_qsys:readdata -> mm_interconnect_1:sysid_qsys_control_slave_readdata
	wire    [0:0] mm_interconnect_1_sysid_qsys_control_slave_address;        // mm_interconnect_1:sysid_qsys_control_slave_address -> sysid_qsys:address
	wire   [31:0] mm_interconnect_1_temp_0_s1_readdata;                      // temp_0:readdata -> mm_interconnect_1:temp_0_s1_readdata
	wire    [1:0] mm_interconnect_1_temp_0_s1_address;                       // mm_interconnect_1:temp_0_s1_address -> temp_0:address
	wire   [31:0] mm_interconnect_1_temp_1_s1_readdata;                      // temp_1:readdata -> mm_interconnect_1:temp_1_s1_readdata
	wire    [1:0] mm_interconnect_1_temp_1_s1_address;                       // mm_interconnect_1:temp_1_s1_address -> temp_1:address
	wire   [31:0] mm_interconnect_1_flags_in_s1_readdata;                    // flags_in:readdata -> mm_interconnect_1:flags_in_s1_readdata
	wire    [1:0] mm_interconnect_1_flags_in_s1_address;                     // mm_interconnect_1:flags_in_s1_address -> flags_in:address
	wire          mm_interconnect_1_flags_out_s1_chipselect;                 // mm_interconnect_1:flags_out_s1_chipselect -> flags_out:chipselect
	wire   [31:0] mm_interconnect_1_flags_out_s1_readdata;                   // flags_out:readdata -> mm_interconnect_1:flags_out_s1_readdata
	wire    [1:0] mm_interconnect_1_flags_out_s1_address;                    // mm_interconnect_1:flags_out_s1_address -> flags_out:address
	wire          mm_interconnect_1_flags_out_s1_write;                      // mm_interconnect_1:flags_out_s1_write -> flags_out:write_n
	wire   [31:0] mm_interconnect_1_flags_out_s1_writedata;                  // mm_interconnect_1:flags_out_s1_writedata -> flags_out:writedata
	wire   [31:0] mm_interconnect_1_temp_2_s1_readdata;                      // temp_2:readdata -> mm_interconnect_1:temp_2_s1_readdata
	wire    [1:0] mm_interconnect_1_temp_2_s1_address;                       // mm_interconnect_1:temp_2_s1_address -> temp_2:address
	wire          mm_interconnect_1_command_type_s1_chipselect;              // mm_interconnect_1:command_type_s1_chipselect -> command_type:chipselect
	wire   [31:0] mm_interconnect_1_command_type_s1_readdata;                // command_type:readdata -> mm_interconnect_1:command_type_s1_readdata
	wire    [1:0] mm_interconnect_1_command_type_s1_address;                 // mm_interconnect_1:command_type_s1_address -> command_type:address
	wire          mm_interconnect_1_command_type_s1_write;                   // mm_interconnect_1:command_type_s1_write -> command_type:write_n
	wire   [31:0] mm_interconnect_1_command_type_s1_writedata;               // mm_interconnect_1:command_type_s1_writedata -> command_type:writedata
	wire          mm_interconnect_1_command_x_s1_chipselect;                 // mm_interconnect_1:command_x_s1_chipselect -> command_x:chipselect
	wire   [31:0] mm_interconnect_1_command_x_s1_readdata;                   // command_x:readdata -> mm_interconnect_1:command_x_s1_readdata
	wire    [1:0] mm_interconnect_1_command_x_s1_address;                    // mm_interconnect_1:command_x_s1_address -> command_x:address
	wire          mm_interconnect_1_command_x_s1_write;                      // mm_interconnect_1:command_x_s1_write -> command_x:write_n
	wire   [31:0] mm_interconnect_1_command_x_s1_writedata;                  // mm_interconnect_1:command_x_s1_writedata -> command_x:writedata
	wire          mm_interconnect_1_command_y_s1_chipselect;                 // mm_interconnect_1:command_y_s1_chipselect -> command_y:chipselect
	wire   [31:0] mm_interconnect_1_command_y_s1_readdata;                   // command_y:readdata -> mm_interconnect_1:command_y_s1_readdata
	wire    [1:0] mm_interconnect_1_command_y_s1_address;                    // mm_interconnect_1:command_y_s1_address -> command_y:address
	wire          mm_interconnect_1_command_y_s1_write;                      // mm_interconnect_1:command_y_s1_write -> command_y:write_n
	wire   [31:0] mm_interconnect_1_command_y_s1_writedata;                  // mm_interconnect_1:command_y_s1_writedata -> command_y:writedata
	wire          mm_interconnect_1_command_z_s1_chipselect;                 // mm_interconnect_1:command_z_s1_chipselect -> command_z:chipselect
	wire   [31:0] mm_interconnect_1_command_z_s1_readdata;                   // command_z:readdata -> mm_interconnect_1:command_z_s1_readdata
	wire    [1:0] mm_interconnect_1_command_z_s1_address;                    // mm_interconnect_1:command_z_s1_address -> command_z:address
	wire          mm_interconnect_1_command_z_s1_write;                      // mm_interconnect_1:command_z_s1_write -> command_z:write_n
	wire   [31:0] mm_interconnect_1_command_z_s1_writedata;                  // mm_interconnect_1:command_z_s1_writedata -> command_z:writedata
	wire          mm_interconnect_1_command_e0_s1_chipselect;                // mm_interconnect_1:command_e0_s1_chipselect -> command_e0:chipselect
	wire   [31:0] mm_interconnect_1_command_e0_s1_readdata;                  // command_e0:readdata -> mm_interconnect_1:command_e0_s1_readdata
	wire    [1:0] mm_interconnect_1_command_e0_s1_address;                   // mm_interconnect_1:command_e0_s1_address -> command_e0:address
	wire          mm_interconnect_1_command_e0_s1_write;                     // mm_interconnect_1:command_e0_s1_write -> command_e0:write_n
	wire   [31:0] mm_interconnect_1_command_e0_s1_writedata;                 // mm_interconnect_1:command_e0_s1_writedata -> command_e0:writedata
	wire          mm_interconnect_1_command_e1_s1_chipselect;                // mm_interconnect_1:command_e1_s1_chipselect -> command_e1:chipselect
	wire   [31:0] mm_interconnect_1_command_e1_s1_readdata;                  // command_e1:readdata -> mm_interconnect_1:command_e1_s1_readdata
	wire    [1:0] mm_interconnect_1_command_e1_s1_address;                   // mm_interconnect_1:command_e1_s1_address -> command_e1:address
	wire          mm_interconnect_1_command_e1_s1_write;                     // mm_interconnect_1:command_e1_s1_write -> command_e1:write_n
	wire   [31:0] mm_interconnect_1_command_e1_s1_writedata;                 // mm_interconnect_1:command_e1_s1_writedata -> command_e1:writedata
	wire          mm_interconnect_1_command_f_x_s1_chipselect;               // mm_interconnect_1:command_f_x_s1_chipselect -> command_f_x:chipselect
	wire   [31:0] mm_interconnect_1_command_f_x_s1_readdata;                 // command_f_x:readdata -> mm_interconnect_1:command_f_x_s1_readdata
	wire    [1:0] mm_interconnect_1_command_f_x_s1_address;                  // mm_interconnect_1:command_f_x_s1_address -> command_f_x:address
	wire          mm_interconnect_1_command_f_x_s1_write;                    // mm_interconnect_1:command_f_x_s1_write -> command_f_x:write_n
	wire   [31:0] mm_interconnect_1_command_f_x_s1_writedata;                // mm_interconnect_1:command_f_x_s1_writedata -> command_f_x:writedata
	wire          mm_interconnect_1_command_t_s1_chipselect;                 // mm_interconnect_1:command_t_s1_chipselect -> command_t:chipselect
	wire   [31:0] mm_interconnect_1_command_t_s1_readdata;                   // command_t:readdata -> mm_interconnect_1:command_t_s1_readdata
	wire    [1:0] mm_interconnect_1_command_t_s1_address;                    // mm_interconnect_1:command_t_s1_address -> command_t:address
	wire          mm_interconnect_1_command_t_s1_write;                      // mm_interconnect_1:command_t_s1_write -> command_t:write_n
	wire   [31:0] mm_interconnect_1_command_t_s1_writedata;                  // mm_interconnect_1:command_t_s1_writedata -> command_t:writedata
	wire          mm_interconnect_1_command_dt_s1_chipselect;                // mm_interconnect_1:command_dt_s1_chipselect -> command_dt:chipselect
	wire   [31:0] mm_interconnect_1_command_dt_s1_readdata;                  // command_dt:readdata -> mm_interconnect_1:command_dt_s1_readdata
	wire    [1:0] mm_interconnect_1_command_dt_s1_address;                   // mm_interconnect_1:command_dt_s1_address -> command_dt:address
	wire          mm_interconnect_1_command_dt_s1_write;                     // mm_interconnect_1:command_dt_s1_write -> command_dt:write_n
	wire   [31:0] mm_interconnect_1_command_dt_s1_writedata;                 // mm_interconnect_1:command_dt_s1_writedata -> command_dt:writedata
	wire          mm_interconnect_1_settings_max_speed_x_s1_chipselect;      // mm_interconnect_1:settings_max_speed_x_s1_chipselect -> settings_max_speed_x:chipselect
	wire   [31:0] mm_interconnect_1_settings_max_speed_x_s1_readdata;        // settings_max_speed_x:readdata -> mm_interconnect_1:settings_max_speed_x_s1_readdata
	wire    [1:0] mm_interconnect_1_settings_max_speed_x_s1_address;         // mm_interconnect_1:settings_max_speed_x_s1_address -> settings_max_speed_x:address
	wire          mm_interconnect_1_settings_max_speed_x_s1_write;           // mm_interconnect_1:settings_max_speed_x_s1_write -> settings_max_speed_x:write_n
	wire   [31:0] mm_interconnect_1_settings_max_speed_x_s1_writedata;       // mm_interconnect_1:settings_max_speed_x_s1_writedata -> settings_max_speed_x:writedata
	wire          mm_interconnect_1_settings_max_speed_y_s1_chipselect;      // mm_interconnect_1:settings_max_speed_y_s1_chipselect -> settings_max_speed_y:chipselect
	wire   [31:0] mm_interconnect_1_settings_max_speed_y_s1_readdata;        // settings_max_speed_y:readdata -> mm_interconnect_1:settings_max_speed_y_s1_readdata
	wire    [1:0] mm_interconnect_1_settings_max_speed_y_s1_address;         // mm_interconnect_1:settings_max_speed_y_s1_address -> settings_max_speed_y:address
	wire          mm_interconnect_1_settings_max_speed_y_s1_write;           // mm_interconnect_1:settings_max_speed_y_s1_write -> settings_max_speed_y:write_n
	wire   [31:0] mm_interconnect_1_settings_max_speed_y_s1_writedata;       // mm_interconnect_1:settings_max_speed_y_s1_writedata -> settings_max_speed_y:writedata
	wire          mm_interconnect_1_settings_max_speed_z_s1_chipselect;      // mm_interconnect_1:settings_max_speed_z_s1_chipselect -> settings_max_speed_z:chipselect
	wire   [31:0] mm_interconnect_1_settings_max_speed_z_s1_readdata;        // settings_max_speed_z:readdata -> mm_interconnect_1:settings_max_speed_z_s1_readdata
	wire    [1:0] mm_interconnect_1_settings_max_speed_z_s1_address;         // mm_interconnect_1:settings_max_speed_z_s1_address -> settings_max_speed_z:address
	wire          mm_interconnect_1_settings_max_speed_z_s1_write;           // mm_interconnect_1:settings_max_speed_z_s1_write -> settings_max_speed_z:write_n
	wire   [31:0] mm_interconnect_1_settings_max_speed_z_s1_writedata;       // mm_interconnect_1:settings_max_speed_z_s1_writedata -> settings_max_speed_z:writedata
	wire          mm_interconnect_1_settings_max_speed_e0_s1_chipselect;     // mm_interconnect_1:settings_max_speed_e0_s1_chipselect -> settings_max_speed_e0:chipselect
	wire   [31:0] mm_interconnect_1_settings_max_speed_e0_s1_readdata;       // settings_max_speed_e0:readdata -> mm_interconnect_1:settings_max_speed_e0_s1_readdata
	wire    [1:0] mm_interconnect_1_settings_max_speed_e0_s1_address;        // mm_interconnect_1:settings_max_speed_e0_s1_address -> settings_max_speed_e0:address
	wire          mm_interconnect_1_settings_max_speed_e0_s1_write;          // mm_interconnect_1:settings_max_speed_e0_s1_write -> settings_max_speed_e0:write_n
	wire   [31:0] mm_interconnect_1_settings_max_speed_e0_s1_writedata;      // mm_interconnect_1:settings_max_speed_e0_s1_writedata -> settings_max_speed_e0:writedata
	wire          mm_interconnect_1_settings_max_speed_e1_s1_chipselect;     // mm_interconnect_1:settings_max_speed_e1_s1_chipselect -> settings_max_speed_e1:chipselect
	wire   [31:0] mm_interconnect_1_settings_max_speed_e1_s1_readdata;       // settings_max_speed_e1:readdata -> mm_interconnect_1:settings_max_speed_e1_s1_readdata
	wire    [1:0] mm_interconnect_1_settings_max_speed_e1_s1_address;        // mm_interconnect_1:settings_max_speed_e1_s1_address -> settings_max_speed_e1:address
	wire          mm_interconnect_1_settings_max_speed_e1_s1_write;          // mm_interconnect_1:settings_max_speed_e1_s1_write -> settings_max_speed_e1:write_n
	wire   [31:0] mm_interconnect_1_settings_max_speed_e1_s1_writedata;      // mm_interconnect_1:settings_max_speed_e1_s1_writedata -> settings_max_speed_e1:writedata
	wire          mm_interconnect_1_settings_acceleration_x_s1_chipselect;   // mm_interconnect_1:settings_acceleration_x_s1_chipselect -> settings_acceleration_x:chipselect
	wire   [31:0] mm_interconnect_1_settings_acceleration_x_s1_readdata;     // settings_acceleration_x:readdata -> mm_interconnect_1:settings_acceleration_x_s1_readdata
	wire    [1:0] mm_interconnect_1_settings_acceleration_x_s1_address;      // mm_interconnect_1:settings_acceleration_x_s1_address -> settings_acceleration_x:address
	wire          mm_interconnect_1_settings_acceleration_x_s1_write;        // mm_interconnect_1:settings_acceleration_x_s1_write -> settings_acceleration_x:write_n
	wire   [31:0] mm_interconnect_1_settings_acceleration_x_s1_writedata;    // mm_interconnect_1:settings_acceleration_x_s1_writedata -> settings_acceleration_x:writedata
	wire          mm_interconnect_1_settings_acceleration_y_s1_chipselect;   // mm_interconnect_1:settings_acceleration_y_s1_chipselect -> settings_acceleration_y:chipselect
	wire   [31:0] mm_interconnect_1_settings_acceleration_y_s1_readdata;     // settings_acceleration_y:readdata -> mm_interconnect_1:settings_acceleration_y_s1_readdata
	wire    [1:0] mm_interconnect_1_settings_acceleration_y_s1_address;      // mm_interconnect_1:settings_acceleration_y_s1_address -> settings_acceleration_y:address
	wire          mm_interconnect_1_settings_acceleration_y_s1_write;        // mm_interconnect_1:settings_acceleration_y_s1_write -> settings_acceleration_y:write_n
	wire   [31:0] mm_interconnect_1_settings_acceleration_y_s1_writedata;    // mm_interconnect_1:settings_acceleration_y_s1_writedata -> settings_acceleration_y:writedata
	wire          mm_interconnect_1_settings_acceleration_e1_s1_chipselect;  // mm_interconnect_1:settings_acceleration_e1_s1_chipselect -> settings_acceleration_e1:chipselect
	wire   [31:0] mm_interconnect_1_settings_acceleration_e1_s1_readdata;    // settings_acceleration_e1:readdata -> mm_interconnect_1:settings_acceleration_e1_s1_readdata
	wire    [1:0] mm_interconnect_1_settings_acceleration_e1_s1_address;     // mm_interconnect_1:settings_acceleration_e1_s1_address -> settings_acceleration_e1:address
	wire          mm_interconnect_1_settings_acceleration_e1_s1_write;       // mm_interconnect_1:settings_acceleration_e1_s1_write -> settings_acceleration_e1:write_n
	wire   [31:0] mm_interconnect_1_settings_acceleration_e1_s1_writedata;   // mm_interconnect_1:settings_acceleration_e1_s1_writedata -> settings_acceleration_e1:writedata
	wire          mm_interconnect_1_settings_acceleration_e0_s1_chipselect;  // mm_interconnect_1:settings_acceleration_e0_s1_chipselect -> settings_acceleration_e0:chipselect
	wire   [31:0] mm_interconnect_1_settings_acceleration_e0_s1_readdata;    // settings_acceleration_e0:readdata -> mm_interconnect_1:settings_acceleration_e0_s1_readdata
	wire    [1:0] mm_interconnect_1_settings_acceleration_e0_s1_address;     // mm_interconnect_1:settings_acceleration_e0_s1_address -> settings_acceleration_e0:address
	wire          mm_interconnect_1_settings_acceleration_e0_s1_write;       // mm_interconnect_1:settings_acceleration_e0_s1_write -> settings_acceleration_e0:write_n
	wire   [31:0] mm_interconnect_1_settings_acceleration_e0_s1_writedata;   // mm_interconnect_1:settings_acceleration_e0_s1_writedata -> settings_acceleration_e0:writedata
	wire          mm_interconnect_1_settings_acceleration_z_s1_chipselect;   // mm_interconnect_1:settings_acceleration_z_s1_chipselect -> settings_acceleration_z:chipselect
	wire   [31:0] mm_interconnect_1_settings_acceleration_z_s1_readdata;     // settings_acceleration_z:readdata -> mm_interconnect_1:settings_acceleration_z_s1_readdata
	wire    [1:0] mm_interconnect_1_settings_acceleration_z_s1_address;      // mm_interconnect_1:settings_acceleration_z_s1_address -> settings_acceleration_z:address
	wire          mm_interconnect_1_settings_acceleration_z_s1_write;        // mm_interconnect_1:settings_acceleration_z_s1_write -> settings_acceleration_z:write_n
	wire   [31:0] mm_interconnect_1_settings_acceleration_z_s1_writedata;    // mm_interconnect_1:settings_acceleration_z_s1_writedata -> settings_acceleration_z:writedata
	wire          mm_interconnect_1_settings_jerk_x_s1_chipselect;           // mm_interconnect_1:settings_jerk_x_s1_chipselect -> settings_jerk_x:chipselect
	wire   [31:0] mm_interconnect_1_settings_jerk_x_s1_readdata;             // settings_jerk_x:readdata -> mm_interconnect_1:settings_jerk_x_s1_readdata
	wire    [1:0] mm_interconnect_1_settings_jerk_x_s1_address;              // mm_interconnect_1:settings_jerk_x_s1_address -> settings_jerk_x:address
	wire          mm_interconnect_1_settings_jerk_x_s1_write;                // mm_interconnect_1:settings_jerk_x_s1_write -> settings_jerk_x:write_n
	wire   [31:0] mm_interconnect_1_settings_jerk_x_s1_writedata;            // mm_interconnect_1:settings_jerk_x_s1_writedata -> settings_jerk_x:writedata
	wire          mm_interconnect_1_settings_jerk_y_s1_chipselect;           // mm_interconnect_1:settings_jerk_y_s1_chipselect -> settings_jerk_y:chipselect
	wire   [31:0] mm_interconnect_1_settings_jerk_y_s1_readdata;             // settings_jerk_y:readdata -> mm_interconnect_1:settings_jerk_y_s1_readdata
	wire    [1:0] mm_interconnect_1_settings_jerk_y_s1_address;              // mm_interconnect_1:settings_jerk_y_s1_address -> settings_jerk_y:address
	wire          mm_interconnect_1_settings_jerk_y_s1_write;                // mm_interconnect_1:settings_jerk_y_s1_write -> settings_jerk_y:write_n
	wire   [31:0] mm_interconnect_1_settings_jerk_y_s1_writedata;            // mm_interconnect_1:settings_jerk_y_s1_writedata -> settings_jerk_y:writedata
	wire          mm_interconnect_1_settings_jerk_z_s1_chipselect;           // mm_interconnect_1:settings_jerk_z_s1_chipselect -> settings_jerk_z:chipselect
	wire   [31:0] mm_interconnect_1_settings_jerk_z_s1_readdata;             // settings_jerk_z:readdata -> mm_interconnect_1:settings_jerk_z_s1_readdata
	wire    [1:0] mm_interconnect_1_settings_jerk_z_s1_address;              // mm_interconnect_1:settings_jerk_z_s1_address -> settings_jerk_z:address
	wire          mm_interconnect_1_settings_jerk_z_s1_write;                // mm_interconnect_1:settings_jerk_z_s1_write -> settings_jerk_z:write_n
	wire   [31:0] mm_interconnect_1_settings_jerk_z_s1_writedata;            // mm_interconnect_1:settings_jerk_z_s1_writedata -> settings_jerk_z:writedata
	wire          mm_interconnect_1_settings_jerk_e0_s1_chipselect;          // mm_interconnect_1:settings_jerk_e0_s1_chipselect -> settings_jerk_e0:chipselect
	wire   [31:0] mm_interconnect_1_settings_jerk_e0_s1_readdata;            // settings_jerk_e0:readdata -> mm_interconnect_1:settings_jerk_e0_s1_readdata
	wire    [1:0] mm_interconnect_1_settings_jerk_e0_s1_address;             // mm_interconnect_1:settings_jerk_e0_s1_address -> settings_jerk_e0:address
	wire          mm_interconnect_1_settings_jerk_e0_s1_write;               // mm_interconnect_1:settings_jerk_e0_s1_write -> settings_jerk_e0:write_n
	wire   [31:0] mm_interconnect_1_settings_jerk_e0_s1_writedata;           // mm_interconnect_1:settings_jerk_e0_s1_writedata -> settings_jerk_e0:writedata
	wire          mm_interconnect_1_settings_jerk_e1_s1_chipselect;          // mm_interconnect_1:settings_jerk_e1_s1_chipselect -> settings_jerk_e1:chipselect
	wire   [31:0] mm_interconnect_1_settings_jerk_e1_s1_readdata;            // settings_jerk_e1:readdata -> mm_interconnect_1:settings_jerk_e1_s1_readdata
	wire    [1:0] mm_interconnect_1_settings_jerk_e1_s1_address;             // mm_interconnect_1:settings_jerk_e1_s1_address -> settings_jerk_e1:address
	wire          mm_interconnect_1_settings_jerk_e1_s1_write;               // mm_interconnect_1:settings_jerk_e1_s1_write -> settings_jerk_e1:write_n
	wire   [31:0] mm_interconnect_1_settings_jerk_e1_s1_writedata;           // mm_interconnect_1:settings_jerk_e1_s1_writedata -> settings_jerk_e1:writedata
	wire          mm_interconnect_1_settings_max_temp_e0_s1_chipselect;      // mm_interconnect_1:settings_max_temp_e0_s1_chipselect -> settings_max_temp_e0:chipselect
	wire   [31:0] mm_interconnect_1_settings_max_temp_e0_s1_readdata;        // settings_max_temp_e0:readdata -> mm_interconnect_1:settings_max_temp_e0_s1_readdata
	wire    [1:0] mm_interconnect_1_settings_max_temp_e0_s1_address;         // mm_interconnect_1:settings_max_temp_e0_s1_address -> settings_max_temp_e0:address
	wire          mm_interconnect_1_settings_max_temp_e0_s1_write;           // mm_interconnect_1:settings_max_temp_e0_s1_write -> settings_max_temp_e0:write_n
	wire   [31:0] mm_interconnect_1_settings_max_temp_e0_s1_writedata;       // mm_interconnect_1:settings_max_temp_e0_s1_writedata -> settings_max_temp_e0:writedata
	wire          mm_interconnect_1_settings_max_temp_e1_s1_chipselect;      // mm_interconnect_1:settings_max_temp_e1_s1_chipselect -> settings_max_temp_e1:chipselect
	wire   [31:0] mm_interconnect_1_settings_max_temp_e1_s1_readdata;        // settings_max_temp_e1:readdata -> mm_interconnect_1:settings_max_temp_e1_s1_readdata
	wire    [1:0] mm_interconnect_1_settings_max_temp_e1_s1_address;         // mm_interconnect_1:settings_max_temp_e1_s1_address -> settings_max_temp_e1:address
	wire          mm_interconnect_1_settings_max_temp_e1_s1_write;           // mm_interconnect_1:settings_max_temp_e1_s1_write -> settings_max_temp_e1:write_n
	wire   [31:0] mm_interconnect_1_settings_max_temp_e1_s1_writedata;       // mm_interconnect_1:settings_max_temp_e1_s1_writedata -> settings_max_temp_e1:writedata
	wire          mm_interconnect_1_settings_max_temp_bed_s1_chipselect;     // mm_interconnect_1:settings_max_temp_bed_s1_chipselect -> settings_max_temp_bed:chipselect
	wire   [31:0] mm_interconnect_1_settings_max_temp_bed_s1_readdata;       // settings_max_temp_bed:readdata -> mm_interconnect_1:settings_max_temp_bed_s1_readdata
	wire    [1:0] mm_interconnect_1_settings_max_temp_bed_s1_address;        // mm_interconnect_1:settings_max_temp_bed_s1_address -> settings_max_temp_bed:address
	wire          mm_interconnect_1_settings_max_temp_bed_s1_write;          // mm_interconnect_1:settings_max_temp_bed_s1_write -> settings_max_temp_bed:write_n
	wire   [31:0] mm_interconnect_1_settings_max_temp_bed_s1_writedata;      // mm_interconnect_1:settings_max_temp_bed_s1_writedata -> settings_max_temp_bed:writedata
	wire   [31:0] mm_interconnect_1_position_x_s1_readdata;                  // position_x:readdata -> mm_interconnect_1:position_x_s1_readdata
	wire    [1:0] mm_interconnect_1_position_x_s1_address;                   // mm_interconnect_1:position_x_s1_address -> position_x:address
	wire   [31:0] mm_interconnect_1_position_y_s1_readdata;                  // position_y:readdata -> mm_interconnect_1:position_y_s1_readdata
	wire    [1:0] mm_interconnect_1_position_y_s1_address;                   // mm_interconnect_1:position_y_s1_address -> position_y:address
	wire   [31:0] mm_interconnect_1_position_z_s1_readdata;                  // position_z:readdata -> mm_interconnect_1:position_z_s1_readdata
	wire    [1:0] mm_interconnect_1_position_z_s1_address;                   // mm_interconnect_1:position_z_s1_address -> position_z:address
	wire   [31:0] mm_interconnect_1_position_e0_s1_readdata;                 // position_e0:readdata -> mm_interconnect_1:position_e0_s1_readdata
	wire    [1:0] mm_interconnect_1_position_e0_s1_address;                  // mm_interconnect_1:position_e0_s1_address -> position_e0:address
	wire   [31:0] mm_interconnect_1_position_e1_s1_readdata;                 // position_e1:readdata -> mm_interconnect_1:position_e1_s1_readdata
	wire    [1:0] mm_interconnect_1_position_e1_s1_address;                  // mm_interconnect_1:position_e1_s1_address -> position_e1:address
	wire          mm_interconnect_1_command_f_y_s1_chipselect;               // mm_interconnect_1:command_f_y_s1_chipselect -> command_f_y:chipselect
	wire   [31:0] mm_interconnect_1_command_f_y_s1_readdata;                 // command_f_y:readdata -> mm_interconnect_1:command_f_y_s1_readdata
	wire    [1:0] mm_interconnect_1_command_f_y_s1_address;                  // mm_interconnect_1:command_f_y_s1_address -> command_f_y:address
	wire          mm_interconnect_1_command_f_y_s1_write;                    // mm_interconnect_1:command_f_y_s1_write -> command_f_y:write_n
	wire   [31:0] mm_interconnect_1_command_f_y_s1_writedata;                // mm_interconnect_1:command_f_y_s1_writedata -> command_f_y:writedata
	wire          mm_interconnect_1_command_f_z_s1_chipselect;               // mm_interconnect_1:command_f_z_s1_chipselect -> command_f_z:chipselect
	wire   [31:0] mm_interconnect_1_command_f_z_s1_readdata;                 // command_f_z:readdata -> mm_interconnect_1:command_f_z_s1_readdata
	wire    [1:0] mm_interconnect_1_command_f_z_s1_address;                  // mm_interconnect_1:command_f_z_s1_address -> command_f_z:address
	wire          mm_interconnect_1_command_f_z_s1_write;                    // mm_interconnect_1:command_f_z_s1_write -> command_f_z:write_n
	wire   [31:0] mm_interconnect_1_command_f_z_s1_writedata;                // mm_interconnect_1:command_f_z_s1_writedata -> command_f_z:writedata
	wire          mm_interconnect_1_command_f_e0_s1_chipselect;              // mm_interconnect_1:command_f_e0_s1_chipselect -> command_f_e0:chipselect
	wire   [31:0] mm_interconnect_1_command_f_e0_s1_readdata;                // command_f_e0:readdata -> mm_interconnect_1:command_f_e0_s1_readdata
	wire    [1:0] mm_interconnect_1_command_f_e0_s1_address;                 // mm_interconnect_1:command_f_e0_s1_address -> command_f_e0:address
	wire          mm_interconnect_1_command_f_e0_s1_write;                   // mm_interconnect_1:command_f_e0_s1_write -> command_f_e0:write_n
	wire   [31:0] mm_interconnect_1_command_f_e0_s1_writedata;               // mm_interconnect_1:command_f_e0_s1_writedata -> command_f_e0:writedata
	wire          mm_interconnect_1_command_f_e1_s1_chipselect;              // mm_interconnect_1:command_f_e1_s1_chipselect -> command_f_e1:chipselect
	wire   [31:0] mm_interconnect_1_command_f_e1_s1_readdata;                // command_f_e1:readdata -> mm_interconnect_1:command_f_e1_s1_readdata
	wire    [1:0] mm_interconnect_1_command_f_e1_s1_address;                 // mm_interconnect_1:command_f_e1_s1_address -> command_f_e1:address
	wire          mm_interconnect_1_command_f_e1_s1_write;                   // mm_interconnect_1:command_f_e1_s1_write -> command_f_e1:write_n
	wire   [31:0] mm_interconnect_1_command_f_e1_s1_writedata;               // mm_interconnect_1:command_f_e1_s1_writedata -> command_f_e1:writedata
	wire   [31:0] mm_interconnect_1_params_x_0_s1_readdata;                  // params_x_0:readdata -> mm_interconnect_1:params_x_0_s1_readdata
	wire    [1:0] mm_interconnect_1_params_x_0_s1_address;                   // mm_interconnect_1:params_x_0_s1_address -> params_x_0:address
	wire   [31:0] mm_interconnect_1_params_x_1_s1_readdata;                  // params_x_1:readdata -> mm_interconnect_1:params_x_1_s1_readdata
	wire    [1:0] mm_interconnect_1_params_x_1_s1_address;                   // mm_interconnect_1:params_x_1_s1_address -> params_x_1:address
	wire   [31:0] mm_interconnect_1_params_x_2_s1_readdata;                  // params_x_2:readdata -> mm_interconnect_1:params_x_2_s1_readdata
	wire    [1:0] mm_interconnect_1_params_x_2_s1_address;                   // mm_interconnect_1:params_x_2_s1_address -> params_x_2:address
	wire   [31:0] mm_interconnect_1_params_x_3_s1_readdata;                  // params_x_3:readdata -> mm_interconnect_1:params_x_3_s1_readdata
	wire    [1:0] mm_interconnect_1_params_x_3_s1_address;                   // mm_interconnect_1:params_x_3_s1_address -> params_x_3:address
	wire   [31:0] mm_interconnect_1_params_x_4_s1_readdata;                  // params_x_4:readdata -> mm_interconnect_1:params_x_4_s1_readdata
	wire    [1:0] mm_interconnect_1_params_x_4_s1_address;                   // mm_interconnect_1:params_x_4_s1_address -> params_x_4:address
	wire   [31:0] mm_interconnect_1_params_y_0_s1_readdata;                  // params_y_0:readdata -> mm_interconnect_1:params_y_0_s1_readdata
	wire    [1:0] mm_interconnect_1_params_y_0_s1_address;                   // mm_interconnect_1:params_y_0_s1_address -> params_y_0:address
	wire   [31:0] mm_interconnect_1_params_y_1_s1_readdata;                  // params_y_1:readdata -> mm_interconnect_1:params_y_1_s1_readdata
	wire    [1:0] mm_interconnect_1_params_y_1_s1_address;                   // mm_interconnect_1:params_y_1_s1_address -> params_y_1:address
	wire   [31:0] mm_interconnect_1_params_y_2_s1_readdata;                  // params_y_2:readdata -> mm_interconnect_1:params_y_2_s1_readdata
	wire    [1:0] mm_interconnect_1_params_y_2_s1_address;                   // mm_interconnect_1:params_y_2_s1_address -> params_y_2:address
	wire   [31:0] mm_interconnect_1_params_y_3_s1_readdata;                  // params_y_3:readdata -> mm_interconnect_1:params_y_3_s1_readdata
	wire    [1:0] mm_interconnect_1_params_y_3_s1_address;                   // mm_interconnect_1:params_y_3_s1_address -> params_y_3:address
	wire   [31:0] mm_interconnect_1_params_y_4_s1_readdata;                  // params_y_4:readdata -> mm_interconnect_1:params_y_4_s1_readdata
	wire    [1:0] mm_interconnect_1_params_y_4_s1_address;                   // mm_interconnect_1:params_y_4_s1_address -> params_y_4:address
	wire   [31:0] mm_interconnect_1_params_z_0_s1_readdata;                  // params_z_0:readdata -> mm_interconnect_1:params_z_0_s1_readdata
	wire    [1:0] mm_interconnect_1_params_z_0_s1_address;                   // mm_interconnect_1:params_z_0_s1_address -> params_z_0:address
	wire   [31:0] mm_interconnect_1_params_z_1_s1_readdata;                  // params_z_1:readdata -> mm_interconnect_1:params_z_1_s1_readdata
	wire    [1:0] mm_interconnect_1_params_z_1_s1_address;                   // mm_interconnect_1:params_z_1_s1_address -> params_z_1:address
	wire   [31:0] mm_interconnect_1_params_z_2_s1_readdata;                  // params_z_2:readdata -> mm_interconnect_1:params_z_2_s1_readdata
	wire    [1:0] mm_interconnect_1_params_z_2_s1_address;                   // mm_interconnect_1:params_z_2_s1_address -> params_z_2:address
	wire   [31:0] mm_interconnect_1_params_z_3_s1_readdata;                  // params_z_3:readdata -> mm_interconnect_1:params_z_3_s1_readdata
	wire    [1:0] mm_interconnect_1_params_z_3_s1_address;                   // mm_interconnect_1:params_z_3_s1_address -> params_z_3:address
	wire   [31:0] mm_interconnect_1_params_z_4_s1_readdata;                  // params_z_4:readdata -> mm_interconnect_1:params_z_4_s1_readdata
	wire    [1:0] mm_interconnect_1_params_z_4_s1_address;                   // mm_interconnect_1:params_z_4_s1_address -> params_z_4:address
	wire   [31:0] mm_interconnect_1_params_e0_0_s1_readdata;                 // params_e0_0:readdata -> mm_interconnect_1:params_e0_0_s1_readdata
	wire    [1:0] mm_interconnect_1_params_e0_0_s1_address;                  // mm_interconnect_1:params_e0_0_s1_address -> params_e0_0:address
	wire   [31:0] mm_interconnect_1_params_e0_1_s1_readdata;                 // params_e0_1:readdata -> mm_interconnect_1:params_e0_1_s1_readdata
	wire    [1:0] mm_interconnect_1_params_e0_1_s1_address;                  // mm_interconnect_1:params_e0_1_s1_address -> params_e0_1:address
	wire   [31:0] mm_interconnect_1_params_e0_2_s1_readdata;                 // params_e0_2:readdata -> mm_interconnect_1:params_e0_2_s1_readdata
	wire    [1:0] mm_interconnect_1_params_e0_2_s1_address;                  // mm_interconnect_1:params_e0_2_s1_address -> params_e0_2:address
	wire   [31:0] mm_interconnect_1_params_e0_3_s1_readdata;                 // params_e0_3:readdata -> mm_interconnect_1:params_e0_3_s1_readdata
	wire    [1:0] mm_interconnect_1_params_e0_3_s1_address;                  // mm_interconnect_1:params_e0_3_s1_address -> params_e0_3:address
	wire   [31:0] mm_interconnect_1_params_e0_4_s1_readdata;                 // params_e0_4:readdata -> mm_interconnect_1:params_e0_4_s1_readdata
	wire    [1:0] mm_interconnect_1_params_e0_4_s1_address;                  // mm_interconnect_1:params_e0_4_s1_address -> params_e0_4:address
	wire   [31:0] mm_interconnect_1_params_e1_0_s1_readdata;                 // params_e1_0:readdata -> mm_interconnect_1:params_e1_0_s1_readdata
	wire    [1:0] mm_interconnect_1_params_e1_0_s1_address;                  // mm_interconnect_1:params_e1_0_s1_address -> params_e1_0:address
	wire   [31:0] mm_interconnect_1_params_e1_4_s1_readdata;                 // params_e1_4:readdata -> mm_interconnect_1:params_e1_4_s1_readdata
	wire    [1:0] mm_interconnect_1_params_e1_4_s1_address;                  // mm_interconnect_1:params_e1_4_s1_address -> params_e1_4:address
	wire   [31:0] mm_interconnect_1_params_e1_3_s1_readdata;                 // params_e1_3:readdata -> mm_interconnect_1:params_e1_3_s1_readdata
	wire    [1:0] mm_interconnect_1_params_e1_3_s1_address;                  // mm_interconnect_1:params_e1_3_s1_address -> params_e1_3:address
	wire   [31:0] mm_interconnect_1_params_e1_2_s1_readdata;                 // params_e1_2:readdata -> mm_interconnect_1:params_e1_2_s1_readdata
	wire    [1:0] mm_interconnect_1_params_e1_2_s1_address;                  // mm_interconnect_1:params_e1_2_s1_address -> params_e1_2:address
	wire   [31:0] mm_interconnect_1_params_e1_1_s1_readdata;                 // params_e1_1:readdata -> mm_interconnect_1:params_e1_1_s1_readdata
	wire    [1:0] mm_interconnect_1_params_e1_1_s1_address;                  // mm_interconnect_1:params_e1_1_s1_address -> params_e1_1:address
	wire   [31:0] mm_interconnect_1_timing_x_0_s1_readdata;                  // timing_x_0:readdata -> mm_interconnect_1:timing_x_0_s1_readdata
	wire    [1:0] mm_interconnect_1_timing_x_0_s1_address;                   // mm_interconnect_1:timing_x_0_s1_address -> timing_x_0:address
	wire   [31:0] mm_interconnect_1_timing_x_1_s1_readdata;                  // timing_x_1:readdata -> mm_interconnect_1:timing_x_1_s1_readdata
	wire    [1:0] mm_interconnect_1_timing_x_1_s1_address;                   // mm_interconnect_1:timing_x_1_s1_address -> timing_x_1:address
	wire   [31:0] mm_interconnect_1_timing_x_2_s1_readdata;                  // timing_x_2:readdata -> mm_interconnect_1:timing_x_2_s1_readdata
	wire    [1:0] mm_interconnect_1_timing_x_2_s1_address;                   // mm_interconnect_1:timing_x_2_s1_address -> timing_x_2:address
	wire   [31:0] mm_interconnect_1_timing_x_3_s1_readdata;                  // timing_x_3:readdata -> mm_interconnect_1:timing_x_3_s1_readdata
	wire    [1:0] mm_interconnect_1_timing_x_3_s1_address;                   // mm_interconnect_1:timing_x_3_s1_address -> timing_x_3:address
	wire   [31:0] mm_interconnect_1_timing_y_0_s1_readdata;                  // timing_y_0:readdata -> mm_interconnect_1:timing_y_0_s1_readdata
	wire    [1:0] mm_interconnect_1_timing_y_0_s1_address;                   // mm_interconnect_1:timing_y_0_s1_address -> timing_y_0:address
	wire   [31:0] mm_interconnect_1_timing_y_1_s1_readdata;                  // timing_y_1:readdata -> mm_interconnect_1:timing_y_1_s1_readdata
	wire    [1:0] mm_interconnect_1_timing_y_1_s1_address;                   // mm_interconnect_1:timing_y_1_s1_address -> timing_y_1:address
	wire   [31:0] mm_interconnect_1_timing_y_2_s1_readdata;                  // timing_y_2:readdata -> mm_interconnect_1:timing_y_2_s1_readdata
	wire    [1:0] mm_interconnect_1_timing_y_2_s1_address;                   // mm_interconnect_1:timing_y_2_s1_address -> timing_y_2:address
	wire   [31:0] mm_interconnect_1_timing_y_3_s1_readdata;                  // timing_y_3:readdata -> mm_interconnect_1:timing_y_3_s1_readdata
	wire    [1:0] mm_interconnect_1_timing_y_3_s1_address;                   // mm_interconnect_1:timing_y_3_s1_address -> timing_y_3:address
	wire   [31:0] mm_interconnect_1_timing_z_0_s1_readdata;                  // timing_z_0:readdata -> mm_interconnect_1:timing_z_0_s1_readdata
	wire    [1:0] mm_interconnect_1_timing_z_0_s1_address;                   // mm_interconnect_1:timing_z_0_s1_address -> timing_z_0:address
	wire   [31:0] mm_interconnect_1_timing_z_1_s1_readdata;                  // timing_z_1:readdata -> mm_interconnect_1:timing_z_1_s1_readdata
	wire    [1:0] mm_interconnect_1_timing_z_1_s1_address;                   // mm_interconnect_1:timing_z_1_s1_address -> timing_z_1:address
	wire   [31:0] mm_interconnect_1_timing_z_2_s1_readdata;                  // timing_z_2:readdata -> mm_interconnect_1:timing_z_2_s1_readdata
	wire    [1:0] mm_interconnect_1_timing_z_2_s1_address;                   // mm_interconnect_1:timing_z_2_s1_address -> timing_z_2:address
	wire   [31:0] mm_interconnect_1_timing_z_3_s1_readdata;                  // timing_z_3:readdata -> mm_interconnect_1:timing_z_3_s1_readdata
	wire    [1:0] mm_interconnect_1_timing_z_3_s1_address;                   // mm_interconnect_1:timing_z_3_s1_address -> timing_z_3:address
	wire   [31:0] mm_interconnect_1_timing_e0_0_s1_readdata;                 // timing_e0_0:readdata -> mm_interconnect_1:timing_e0_0_s1_readdata
	wire    [1:0] mm_interconnect_1_timing_e0_0_s1_address;                  // mm_interconnect_1:timing_e0_0_s1_address -> timing_e0_0:address
	wire   [31:0] mm_interconnect_1_timing_e0_1_s1_readdata;                 // timing_e0_1:readdata -> mm_interconnect_1:timing_e0_1_s1_readdata
	wire    [1:0] mm_interconnect_1_timing_e0_1_s1_address;                  // mm_interconnect_1:timing_e0_1_s1_address -> timing_e0_1:address
	wire   [31:0] mm_interconnect_1_timing_e0_2_s1_readdata;                 // timing_e0_2:readdata -> mm_interconnect_1:timing_e0_2_s1_readdata
	wire    [1:0] mm_interconnect_1_timing_e0_2_s1_address;                  // mm_interconnect_1:timing_e0_2_s1_address -> timing_e0_2:address
	wire   [31:0] mm_interconnect_1_timing_e0_3_s1_readdata;                 // timing_e0_3:readdata -> mm_interconnect_1:timing_e0_3_s1_readdata
	wire    [1:0] mm_interconnect_1_timing_e0_3_s1_address;                  // mm_interconnect_1:timing_e0_3_s1_address -> timing_e0_3:address
	wire   [31:0] mm_interconnect_1_timing_e1_0_s1_readdata;                 // timing_e1_0:readdata -> mm_interconnect_1:timing_e1_0_s1_readdata
	wire    [1:0] mm_interconnect_1_timing_e1_0_s1_address;                  // mm_interconnect_1:timing_e1_0_s1_address -> timing_e1_0:address
	wire   [31:0] mm_interconnect_1_timing_e1_1_s1_readdata;                 // timing_e1_1:readdata -> mm_interconnect_1:timing_e1_1_s1_readdata
	wire    [1:0] mm_interconnect_1_timing_e1_1_s1_address;                  // mm_interconnect_1:timing_e1_1_s1_address -> timing_e1_1:address
	wire   [31:0] mm_interconnect_1_timing_e1_2_s1_readdata;                 // timing_e1_2:readdata -> mm_interconnect_1:timing_e1_2_s1_readdata
	wire    [1:0] mm_interconnect_1_timing_e1_2_s1_address;                  // mm_interconnect_1:timing_e1_2_s1_address -> timing_e1_2:address
	wire   [31:0] mm_interconnect_1_timing_e1_3_s1_readdata;                 // timing_e1_3:readdata -> mm_interconnect_1:timing_e1_3_s1_readdata
	wire    [1:0] mm_interconnect_1_timing_e1_3_s1_address;                  // mm_interconnect_1:timing_e1_3_s1_address -> timing_e1_3:address
	wire   [31:0] mm_interconnect_1_new_rparams_x_0_s1_readdata;             // new_rparams_x_0:readdata -> mm_interconnect_1:new_rparams_x_0_s1_readdata
	wire    [1:0] mm_interconnect_1_new_rparams_x_0_s1_address;              // mm_interconnect_1:new_rparams_x_0_s1_address -> new_rparams_x_0:address
	wire   [31:0] mm_interconnect_1_new_rparams_x_1_s1_readdata;             // new_rparams_x_1:readdata -> mm_interconnect_1:new_rparams_x_1_s1_readdata
	wire    [1:0] mm_interconnect_1_new_rparams_x_1_s1_address;              // mm_interconnect_1:new_rparams_x_1_s1_address -> new_rparams_x_1:address
	wire   [31:0] mm_interconnect_1_new_rparams_x_2_s1_readdata;             // new_rparams_x_2:readdata -> mm_interconnect_1:new_rparams_x_2_s1_readdata
	wire    [1:0] mm_interconnect_1_new_rparams_x_2_s1_address;              // mm_interconnect_1:new_rparams_x_2_s1_address -> new_rparams_x_2:address
	wire   [31:0] mm_interconnect_1_new_rparams_x_3_s1_readdata;             // new_rparams_x_3:readdata -> mm_interconnect_1:new_rparams_x_3_s1_readdata
	wire    [1:0] mm_interconnect_1_new_rparams_x_3_s1_address;              // mm_interconnect_1:new_rparams_x_3_s1_address -> new_rparams_x_3:address
	wire   [31:0] mm_interconnect_1_new_rparams_x_4_s1_readdata;             // new_rparams_x_4:readdata -> mm_interconnect_1:new_rparams_x_4_s1_readdata
	wire    [1:0] mm_interconnect_1_new_rparams_x_4_s1_address;              // mm_interconnect_1:new_rparams_x_4_s1_address -> new_rparams_x_4:address
	wire   [31:0] mm_interconnect_1_new_rparams_y_0_s1_readdata;             // new_rparams_y_0:readdata -> mm_interconnect_1:new_rparams_y_0_s1_readdata
	wire    [1:0] mm_interconnect_1_new_rparams_y_0_s1_address;              // mm_interconnect_1:new_rparams_y_0_s1_address -> new_rparams_y_0:address
	wire   [31:0] mm_interconnect_1_new_rparams_y_1_s1_readdata;             // new_rparams_y_1:readdata -> mm_interconnect_1:new_rparams_y_1_s1_readdata
	wire    [1:0] mm_interconnect_1_new_rparams_y_1_s1_address;              // mm_interconnect_1:new_rparams_y_1_s1_address -> new_rparams_y_1:address
	wire   [31:0] mm_interconnect_1_new_rparams_y_2_s1_readdata;             // new_rparams_y_2:readdata -> mm_interconnect_1:new_rparams_y_2_s1_readdata
	wire    [1:0] mm_interconnect_1_new_rparams_y_2_s1_address;              // mm_interconnect_1:new_rparams_y_2_s1_address -> new_rparams_y_2:address
	wire   [31:0] mm_interconnect_1_new_rparams_y_3_s1_readdata;             // new_rparams_y_3:readdata -> mm_interconnect_1:new_rparams_y_3_s1_readdata
	wire    [1:0] mm_interconnect_1_new_rparams_y_3_s1_address;              // mm_interconnect_1:new_rparams_y_3_s1_address -> new_rparams_y_3:address
	wire   [31:0] mm_interconnect_1_new_rparams_y_4_s1_readdata;             // new_rparams_y_4:readdata -> mm_interconnect_1:new_rparams_y_4_s1_readdata
	wire    [1:0] mm_interconnect_1_new_rparams_y_4_s1_address;              // mm_interconnect_1:new_rparams_y_4_s1_address -> new_rparams_y_4:address
	wire   [31:0] mm_interconnect_1_new_rparams_z_0_s1_readdata;             // new_rparams_z_0:readdata -> mm_interconnect_1:new_rparams_z_0_s1_readdata
	wire    [1:0] mm_interconnect_1_new_rparams_z_0_s1_address;              // mm_interconnect_1:new_rparams_z_0_s1_address -> new_rparams_z_0:address
	wire   [31:0] mm_interconnect_1_new_rparams_z_1_s1_readdata;             // new_rparams_z_1:readdata -> mm_interconnect_1:new_rparams_z_1_s1_readdata
	wire    [1:0] mm_interconnect_1_new_rparams_z_1_s1_address;              // mm_interconnect_1:new_rparams_z_1_s1_address -> new_rparams_z_1:address
	wire   [31:0] mm_interconnect_1_new_rparams_z_2_s1_readdata;             // new_rparams_z_2:readdata -> mm_interconnect_1:new_rparams_z_2_s1_readdata
	wire    [1:0] mm_interconnect_1_new_rparams_z_2_s1_address;              // mm_interconnect_1:new_rparams_z_2_s1_address -> new_rparams_z_2:address
	wire   [31:0] mm_interconnect_1_new_rparams_z_3_s1_readdata;             // new_rparams_z_3:readdata -> mm_interconnect_1:new_rparams_z_3_s1_readdata
	wire    [1:0] mm_interconnect_1_new_rparams_z_3_s1_address;              // mm_interconnect_1:new_rparams_z_3_s1_address -> new_rparams_z_3:address
	wire   [31:0] mm_interconnect_1_new_rparams_z_4_s1_readdata;             // new_rparams_z_4:readdata -> mm_interconnect_1:new_rparams_z_4_s1_readdata
	wire    [1:0] mm_interconnect_1_new_rparams_z_4_s1_address;              // mm_interconnect_1:new_rparams_z_4_s1_address -> new_rparams_z_4:address
	wire   [31:0] mm_interconnect_1_new_rparams_e0_0_s1_readdata;            // new_rparams_e0_0:readdata -> mm_interconnect_1:new_rparams_e0_0_s1_readdata
	wire    [1:0] mm_interconnect_1_new_rparams_e0_0_s1_address;             // mm_interconnect_1:new_rparams_e0_0_s1_address -> new_rparams_e0_0:address
	wire   [31:0] mm_interconnect_1_new_rparams_e0_1_s1_readdata;            // new_rparams_e0_1:readdata -> mm_interconnect_1:new_rparams_e0_1_s1_readdata
	wire    [1:0] mm_interconnect_1_new_rparams_e0_1_s1_address;             // mm_interconnect_1:new_rparams_e0_1_s1_address -> new_rparams_e0_1:address
	wire   [31:0] mm_interconnect_1_new_rparams_e0_2_s1_readdata;            // new_rparams_e0_2:readdata -> mm_interconnect_1:new_rparams_e0_2_s1_readdata
	wire    [1:0] mm_interconnect_1_new_rparams_e0_2_s1_address;             // mm_interconnect_1:new_rparams_e0_2_s1_address -> new_rparams_e0_2:address
	wire   [31:0] mm_interconnect_1_new_rparams_e0_3_s1_readdata;            // new_rparams_e0_3:readdata -> mm_interconnect_1:new_rparams_e0_3_s1_readdata
	wire    [1:0] mm_interconnect_1_new_rparams_e0_3_s1_address;             // mm_interconnect_1:new_rparams_e0_3_s1_address -> new_rparams_e0_3:address
	wire   [31:0] mm_interconnect_1_new_rparams_e0_4_s1_readdata;            // new_rparams_e0_4:readdata -> mm_interconnect_1:new_rparams_e0_4_s1_readdata
	wire    [1:0] mm_interconnect_1_new_rparams_e0_4_s1_address;             // mm_interconnect_1:new_rparams_e0_4_s1_address -> new_rparams_e0_4:address
	wire   [31:0] mm_interconnect_1_new_rparams_e1_0_s1_readdata;            // new_rparams_e1_0:readdata -> mm_interconnect_1:new_rparams_e1_0_s1_readdata
	wire    [1:0] mm_interconnect_1_new_rparams_e1_0_s1_address;             // mm_interconnect_1:new_rparams_e1_0_s1_address -> new_rparams_e1_0:address
	wire   [31:0] mm_interconnect_1_new_rparams_e1_1_s1_readdata;            // new_rparams_e1_1:readdata -> mm_interconnect_1:new_rparams_e1_1_s1_readdata
	wire    [1:0] mm_interconnect_1_new_rparams_e1_1_s1_address;             // mm_interconnect_1:new_rparams_e1_1_s1_address -> new_rparams_e1_1:address
	wire   [31:0] mm_interconnect_1_new_rparams_e1_2_s1_readdata;            // new_rparams_e1_2:readdata -> mm_interconnect_1:new_rparams_e1_2_s1_readdata
	wire    [1:0] mm_interconnect_1_new_rparams_e1_2_s1_address;             // mm_interconnect_1:new_rparams_e1_2_s1_address -> new_rparams_e1_2:address
	wire   [31:0] mm_interconnect_1_new_rparams_e1_3_s1_readdata;            // new_rparams_e1_3:readdata -> mm_interconnect_1:new_rparams_e1_3_s1_readdata
	wire    [1:0] mm_interconnect_1_new_rparams_e1_3_s1_address;             // mm_interconnect_1:new_rparams_e1_3_s1_address -> new_rparams_e1_3:address
	wire   [31:0] mm_interconnect_1_new_rparams_e1_4_s1_readdata;            // new_rparams_e1_4:readdata -> mm_interconnect_1:new_rparams_e1_4_s1_readdata
	wire    [1:0] mm_interconnect_1_new_rparams_e1_4_s1_address;             // mm_interconnect_1:new_rparams_e1_4_s1_address -> new_rparams_e1_4:address
	wire   [31:0] mm_interconnect_1_step_x_now_s1_readdata;                  // step_x_now:readdata -> mm_interconnect_1:step_x_now_s1_readdata
	wire    [1:0] mm_interconnect_1_step_x_now_s1_address;                   // mm_interconnect_1:step_x_now_s1_address -> step_x_now:address
	wire   [31:0] mm_interconnect_1_step_y_now_s1_readdata;                  // step_y_now:readdata -> mm_interconnect_1:step_y_now_s1_readdata
	wire    [1:0] mm_interconnect_1_step_y_now_s1_address;                   // mm_interconnect_1:step_y_now_s1_address -> step_y_now:address
	wire   [31:0] mm_interconnect_1_step_z_now_s1_readdata;                  // step_z_now:readdata -> mm_interconnect_1:step_z_now_s1_readdata
	wire    [1:0] mm_interconnect_1_step_z_now_s1_address;                   // mm_interconnect_1:step_z_now_s1_address -> step_z_now:address
	wire   [31:0] mm_interconnect_1_step_e0_now_s1_readdata;                 // step_e0_now:readdata -> mm_interconnect_1:step_e0_now_s1_readdata
	wire    [1:0] mm_interconnect_1_step_e0_now_s1_address;                  // mm_interconnect_1:step_e0_now_s1_address -> step_e0_now:address
	wire   [31:0] mm_interconnect_1_step_e1_now_s1_readdata;                 // step_e1_now:readdata -> mm_interconnect_1:step_e1_now_s1_readdata
	wire    [1:0] mm_interconnect_1_step_e1_now_s1_address;                  // mm_interconnect_1:step_e1_now_s1_address -> step_e1_now:address
	wire   [31:0] mm_interconnect_1_max_params_0_s1_readdata;                // max_params_0:readdata -> mm_interconnect_1:max_params_0_s1_readdata
	wire    [1:0] mm_interconnect_1_max_params_0_s1_address;                 // mm_interconnect_1:max_params_0_s1_address -> max_params_0:address
	wire   [31:0] mm_interconnect_1_max_params_1_s1_readdata;                // max_params_1:readdata -> mm_interconnect_1:max_params_1_s1_readdata
	wire    [1:0] mm_interconnect_1_max_params_1_s1_address;                 // mm_interconnect_1:max_params_1_s1_address -> max_params_1:address
	wire   [31:0] mm_interconnect_1_max_params_2_s1_readdata;                // max_params_2:readdata -> mm_interconnect_1:max_params_2_s1_readdata
	wire    [1:0] mm_interconnect_1_max_params_2_s1_address;                 // mm_interconnect_1:max_params_2_s1_address -> max_params_2:address
	wire   [31:0] mm_interconnect_1_max_params_3_s1_readdata;                // max_params_3:readdata -> mm_interconnect_1:max_params_3_s1_readdata
	wire    [1:0] mm_interconnect_1_max_params_3_s1_address;                 // mm_interconnect_1:max_params_3_s1_address -> max_params_3:address
	wire   [31:0] mm_interconnect_1_max_params_4_s1_readdata;                // max_params_4:readdata -> mm_interconnect_1:max_params_4_s1_readdata
	wire    [1:0] mm_interconnect_1_max_params_4_s1_address;                 // mm_interconnect_1:max_params_4_s1_address -> max_params_4:address
	wire   [31:0] mm_interconnect_1_max_timing_0_s1_readdata;                // max_timing_0:readdata -> mm_interconnect_1:max_timing_0_s1_readdata
	wire    [1:0] mm_interconnect_1_max_timing_0_s1_address;                 // mm_interconnect_1:max_timing_0_s1_address -> max_timing_0:address
	wire   [31:0] mm_interconnect_1_max_timing_3_s1_readdata;                // max_timing_3:readdata -> mm_interconnect_1:max_timing_3_s1_readdata
	wire    [1:0] mm_interconnect_1_max_timing_3_s1_address;                 // mm_interconnect_1:max_timing_3_s1_address -> max_timing_3:address
	wire   [31:0] mm_interconnect_1_max_timing_2_s1_readdata;                // max_timing_2:readdata -> mm_interconnect_1:max_timing_2_s1_readdata
	wire    [1:0] mm_interconnect_1_max_timing_2_s1_address;                 // mm_interconnect_1:max_timing_2_s1_address -> max_timing_2:address
	wire   [31:0] mm_interconnect_1_max_timing_1_s1_readdata;                // max_timing_1:readdata -> mm_interconnect_1:max_timing_1_s1_readdata
	wire    [1:0] mm_interconnect_1_max_timing_1_s1_address;                 // mm_interconnect_1:max_timing_1_s1_address -> max_timing_1:address
	wire   [31:0] hps_only_master_master_readdata;                           // mm_interconnect_2:hps_only_master_master_readdata -> hps_only_master:master_readdata
	wire          hps_only_master_master_waitrequest;                        // mm_interconnect_2:hps_only_master_master_waitrequest -> hps_only_master:master_waitrequest
	wire   [31:0] hps_only_master_master_address;                            // hps_only_master:master_address -> mm_interconnect_2:hps_only_master_master_address
	wire          hps_only_master_master_read;                               // hps_only_master:master_read -> mm_interconnect_2:hps_only_master_master_read
	wire    [3:0] hps_only_master_master_byteenable;                         // hps_only_master:master_byteenable -> mm_interconnect_2:hps_only_master_master_byteenable
	wire          hps_only_master_master_readdatavalid;                      // mm_interconnect_2:hps_only_master_master_readdatavalid -> hps_only_master:master_readdatavalid
	wire          hps_only_master_master_write;                              // hps_only_master:master_write -> mm_interconnect_2:hps_only_master_master_write
	wire   [31:0] hps_only_master_master_writedata;                          // hps_only_master:master_writedata -> mm_interconnect_2:hps_only_master_master_writedata
	wire    [1:0] mm_interconnect_2_hps_0_f2h_axi_slave_awburst;             // mm_interconnect_2:hps_0_f2h_axi_slave_awburst -> hps_0:f2h_AWBURST
	wire    [4:0] mm_interconnect_2_hps_0_f2h_axi_slave_awuser;              // mm_interconnect_2:hps_0_f2h_axi_slave_awuser -> hps_0:f2h_AWUSER
	wire    [3:0] mm_interconnect_2_hps_0_f2h_axi_slave_arlen;               // mm_interconnect_2:hps_0_f2h_axi_slave_arlen -> hps_0:f2h_ARLEN
	wire    [7:0] mm_interconnect_2_hps_0_f2h_axi_slave_wstrb;               // mm_interconnect_2:hps_0_f2h_axi_slave_wstrb -> hps_0:f2h_WSTRB
	wire          mm_interconnect_2_hps_0_f2h_axi_slave_wready;              // hps_0:f2h_WREADY -> mm_interconnect_2:hps_0_f2h_axi_slave_wready
	wire    [7:0] mm_interconnect_2_hps_0_f2h_axi_slave_rid;                 // hps_0:f2h_RID -> mm_interconnect_2:hps_0_f2h_axi_slave_rid
	wire          mm_interconnect_2_hps_0_f2h_axi_slave_rready;              // mm_interconnect_2:hps_0_f2h_axi_slave_rready -> hps_0:f2h_RREADY
	wire    [3:0] mm_interconnect_2_hps_0_f2h_axi_slave_awlen;               // mm_interconnect_2:hps_0_f2h_axi_slave_awlen -> hps_0:f2h_AWLEN
	wire    [7:0] mm_interconnect_2_hps_0_f2h_axi_slave_wid;                 // mm_interconnect_2:hps_0_f2h_axi_slave_wid -> hps_0:f2h_WID
	wire    [3:0] mm_interconnect_2_hps_0_f2h_axi_slave_arcache;             // mm_interconnect_2:hps_0_f2h_axi_slave_arcache -> hps_0:f2h_ARCACHE
	wire          mm_interconnect_2_hps_0_f2h_axi_slave_wvalid;              // mm_interconnect_2:hps_0_f2h_axi_slave_wvalid -> hps_0:f2h_WVALID
	wire   [31:0] mm_interconnect_2_hps_0_f2h_axi_slave_araddr;              // mm_interconnect_2:hps_0_f2h_axi_slave_araddr -> hps_0:f2h_ARADDR
	wire    [2:0] mm_interconnect_2_hps_0_f2h_axi_slave_arprot;              // mm_interconnect_2:hps_0_f2h_axi_slave_arprot -> hps_0:f2h_ARPROT
	wire    [2:0] mm_interconnect_2_hps_0_f2h_axi_slave_awprot;              // mm_interconnect_2:hps_0_f2h_axi_slave_awprot -> hps_0:f2h_AWPROT
	wire   [63:0] mm_interconnect_2_hps_0_f2h_axi_slave_wdata;               // mm_interconnect_2:hps_0_f2h_axi_slave_wdata -> hps_0:f2h_WDATA
	wire          mm_interconnect_2_hps_0_f2h_axi_slave_arvalid;             // mm_interconnect_2:hps_0_f2h_axi_slave_arvalid -> hps_0:f2h_ARVALID
	wire    [3:0] mm_interconnect_2_hps_0_f2h_axi_slave_awcache;             // mm_interconnect_2:hps_0_f2h_axi_slave_awcache -> hps_0:f2h_AWCACHE
	wire    [7:0] mm_interconnect_2_hps_0_f2h_axi_slave_arid;                // mm_interconnect_2:hps_0_f2h_axi_slave_arid -> hps_0:f2h_ARID
	wire    [1:0] mm_interconnect_2_hps_0_f2h_axi_slave_arlock;              // mm_interconnect_2:hps_0_f2h_axi_slave_arlock -> hps_0:f2h_ARLOCK
	wire    [1:0] mm_interconnect_2_hps_0_f2h_axi_slave_awlock;              // mm_interconnect_2:hps_0_f2h_axi_slave_awlock -> hps_0:f2h_AWLOCK
	wire   [31:0] mm_interconnect_2_hps_0_f2h_axi_slave_awaddr;              // mm_interconnect_2:hps_0_f2h_axi_slave_awaddr -> hps_0:f2h_AWADDR
	wire    [1:0] mm_interconnect_2_hps_0_f2h_axi_slave_bresp;               // hps_0:f2h_BRESP -> mm_interconnect_2:hps_0_f2h_axi_slave_bresp
	wire          mm_interconnect_2_hps_0_f2h_axi_slave_arready;             // hps_0:f2h_ARREADY -> mm_interconnect_2:hps_0_f2h_axi_slave_arready
	wire   [63:0] mm_interconnect_2_hps_0_f2h_axi_slave_rdata;               // hps_0:f2h_RDATA -> mm_interconnect_2:hps_0_f2h_axi_slave_rdata
	wire          mm_interconnect_2_hps_0_f2h_axi_slave_awready;             // hps_0:f2h_AWREADY -> mm_interconnect_2:hps_0_f2h_axi_slave_awready
	wire    [1:0] mm_interconnect_2_hps_0_f2h_axi_slave_arburst;             // mm_interconnect_2:hps_0_f2h_axi_slave_arburst -> hps_0:f2h_ARBURST
	wire    [2:0] mm_interconnect_2_hps_0_f2h_axi_slave_arsize;              // mm_interconnect_2:hps_0_f2h_axi_slave_arsize -> hps_0:f2h_ARSIZE
	wire          mm_interconnect_2_hps_0_f2h_axi_slave_bready;              // mm_interconnect_2:hps_0_f2h_axi_slave_bready -> hps_0:f2h_BREADY
	wire          mm_interconnect_2_hps_0_f2h_axi_slave_rlast;               // hps_0:f2h_RLAST -> mm_interconnect_2:hps_0_f2h_axi_slave_rlast
	wire          mm_interconnect_2_hps_0_f2h_axi_slave_wlast;               // mm_interconnect_2:hps_0_f2h_axi_slave_wlast -> hps_0:f2h_WLAST
	wire    [1:0] mm_interconnect_2_hps_0_f2h_axi_slave_rresp;               // hps_0:f2h_RRESP -> mm_interconnect_2:hps_0_f2h_axi_slave_rresp
	wire    [7:0] mm_interconnect_2_hps_0_f2h_axi_slave_awid;                // mm_interconnect_2:hps_0_f2h_axi_slave_awid -> hps_0:f2h_AWID
	wire    [7:0] mm_interconnect_2_hps_0_f2h_axi_slave_bid;                 // hps_0:f2h_BID -> mm_interconnect_2:hps_0_f2h_axi_slave_bid
	wire          mm_interconnect_2_hps_0_f2h_axi_slave_bvalid;              // hps_0:f2h_BVALID -> mm_interconnect_2:hps_0_f2h_axi_slave_bvalid
	wire    [2:0] mm_interconnect_2_hps_0_f2h_axi_slave_awsize;              // mm_interconnect_2:hps_0_f2h_axi_slave_awsize -> hps_0:f2h_AWSIZE
	wire          mm_interconnect_2_hps_0_f2h_axi_slave_awvalid;             // mm_interconnect_2:hps_0_f2h_axi_slave_awvalid -> hps_0:f2h_AWVALID
	wire    [4:0] mm_interconnect_2_hps_0_f2h_axi_slave_aruser;              // mm_interconnect_2:hps_0_f2h_axi_slave_aruser -> hps_0:f2h_ARUSER
	wire          mm_interconnect_2_hps_0_f2h_axi_slave_rvalid;              // hps_0:f2h_RVALID -> mm_interconnect_2:hps_0_f2h_axi_slave_rvalid
	wire   [31:0] f2sdram_only_master_master_readdata;                       // mm_interconnect_3:f2sdram_only_master_master_readdata -> f2sdram_only_master:master_readdata
	wire          f2sdram_only_master_master_waitrequest;                    // mm_interconnect_3:f2sdram_only_master_master_waitrequest -> f2sdram_only_master:master_waitrequest
	wire   [31:0] f2sdram_only_master_master_address;                        // f2sdram_only_master:master_address -> mm_interconnect_3:f2sdram_only_master_master_address
	wire          f2sdram_only_master_master_read;                           // f2sdram_only_master:master_read -> mm_interconnect_3:f2sdram_only_master_master_read
	wire    [3:0] f2sdram_only_master_master_byteenable;                     // f2sdram_only_master:master_byteenable -> mm_interconnect_3:f2sdram_only_master_master_byteenable
	wire          f2sdram_only_master_master_readdatavalid;                  // mm_interconnect_3:f2sdram_only_master_master_readdatavalid -> f2sdram_only_master:master_readdatavalid
	wire          f2sdram_only_master_master_write;                          // f2sdram_only_master:master_write -> mm_interconnect_3:f2sdram_only_master_master_write
	wire   [31:0] f2sdram_only_master_master_writedata;                      // f2sdram_only_master:master_writedata -> mm_interconnect_3:f2sdram_only_master_master_writedata
	wire  [255:0] mm_interconnect_3_hps_0_f2h_sdram0_data_readdata;          // hps_0:f2h_sdram0_READDATA -> mm_interconnect_3:hps_0_f2h_sdram0_data_readdata
	wire          mm_interconnect_3_hps_0_f2h_sdram0_data_waitrequest;       // hps_0:f2h_sdram0_WAITREQUEST -> mm_interconnect_3:hps_0_f2h_sdram0_data_waitrequest
	wire   [26:0] mm_interconnect_3_hps_0_f2h_sdram0_data_address;           // mm_interconnect_3:hps_0_f2h_sdram0_data_address -> hps_0:f2h_sdram0_ADDRESS
	wire          mm_interconnect_3_hps_0_f2h_sdram0_data_read;              // mm_interconnect_3:hps_0_f2h_sdram0_data_read -> hps_0:f2h_sdram0_READ
	wire   [31:0] mm_interconnect_3_hps_0_f2h_sdram0_data_byteenable;        // mm_interconnect_3:hps_0_f2h_sdram0_data_byteenable -> hps_0:f2h_sdram0_BYTEENABLE
	wire          mm_interconnect_3_hps_0_f2h_sdram0_data_readdatavalid;     // hps_0:f2h_sdram0_READDATAVALID -> mm_interconnect_3:hps_0_f2h_sdram0_data_readdatavalid
	wire          mm_interconnect_3_hps_0_f2h_sdram0_data_write;             // mm_interconnect_3:hps_0_f2h_sdram0_data_write -> hps_0:f2h_sdram0_WRITE
	wire  [255:0] mm_interconnect_3_hps_0_f2h_sdram0_data_writedata;         // mm_interconnect_3:hps_0_f2h_sdram0_data_writedata -> hps_0:f2h_sdram0_WRITEDATA
	wire    [7:0] mm_interconnect_3_hps_0_f2h_sdram0_data_burstcount;        // mm_interconnect_3:hps_0_f2h_sdram0_data_burstcount -> hps_0:f2h_sdram0_BURSTCOUNT
	wire    [2:0] ilc_irq_irq;                                               // irq_mapper:sender_irq -> ILC:irq
	wire   [31:0] hps_0_f2h_irq0_irq;                                        // irq_mapper_001:sender_irq -> hps_0:f2h_irq_p0
	wire   [31:0] hps_0_f2h_irq1_irq;                                        // irq_mapper_002:sender_irq -> hps_0:f2h_irq_p1
	wire          irq_mapper_receiver0_irq;                                  // jtag_uart:av_irq -> [irq_mapper:receiver0_irq, irq_mapper_001:receiver0_irq]
	wire          rst_controller_reset_out_reset;                            // rst_controller:reset_out -> [ILC:reset_n, command_dt:reset_n, command_e0:reset_n, command_e1:reset_n, command_f_e0:reset_n, command_f_e1:reset_n, command_f_x:reset_n, command_f_y:reset_n, command_f_z:reset_n, command_t:reset_n, command_type:reset_n, command_x:reset_n, command_y:reset_n, command_z:reset_n, flags_in:reset_n, flags_out:reset_n, irq_mapper:reset, jtag_uart:rst_n, max_params_0:reset_n, max_params_1:reset_n, max_params_2:reset_n, max_params_3:reset_n, max_params_4:reset_n, max_timing_0:reset_n, max_timing_1:reset_n, max_timing_2:reset_n, max_timing_3:reset_n, mm_bridge_0:reset, mm_interconnect_0:mm_bridge_0_reset_reset_bridge_in_reset_reset, mm_interconnect_1:fpga_only_master_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_1:mm_bridge_0_reset_reset_bridge_in_reset_reset, mm_interconnect_2:hps_only_master_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_2:hps_only_master_master_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_3:f2sdram_only_master_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_3:f2sdram_only_master_master_translator_reset_reset_bridge_in_reset_reset, new_rparams_e0_0:reset_n, new_rparams_e0_1:reset_n, new_rparams_e0_2:reset_n, new_rparams_e0_3:reset_n, new_rparams_e0_4:reset_n, new_rparams_e1_0:reset_n, new_rparams_e1_1:reset_n, new_rparams_e1_2:reset_n, new_rparams_e1_3:reset_n, new_rparams_e1_4:reset_n, new_rparams_x_0:reset_n, new_rparams_x_1:reset_n, new_rparams_x_2:reset_n, new_rparams_x_3:reset_n, new_rparams_x_4:reset_n, new_rparams_y_0:reset_n, new_rparams_y_1:reset_n, new_rparams_y_2:reset_n, new_rparams_y_3:reset_n, new_rparams_y_4:reset_n, new_rparams_z_0:reset_n, new_rparams_z_1:reset_n, new_rparams_z_2:reset_n, new_rparams_z_3:reset_n, new_rparams_z_4:reset_n, params_e0_0:reset_n, params_e0_1:reset_n, params_e0_2:reset_n, params_e0_3:reset_n, params_e0_4:reset_n, params_e1_0:reset_n, params_e1_1:reset_n, params_e1_2:reset_n, params_e1_3:reset_n, params_e1_4:reset_n, params_x_0:reset_n, params_x_1:reset_n, params_x_2:reset_n, params_x_3:reset_n, params_x_4:reset_n, params_y_0:reset_n, params_y_1:reset_n, params_y_2:reset_n, params_y_3:reset_n, params_y_4:reset_n, params_z_0:reset_n, params_z_1:reset_n, params_z_2:reset_n, params_z_3:reset_n, params_z_4:reset_n, position_e0:reset_n, position_e1:reset_n, position_x:reset_n, position_y:reset_n, position_z:reset_n, settings_acceleration_e0:reset_n, settings_acceleration_e1:reset_n, settings_acceleration_x:reset_n, settings_acceleration_y:reset_n, settings_acceleration_z:reset_n, settings_jerk_e0:reset_n, settings_jerk_e1:reset_n, settings_jerk_x:reset_n, settings_jerk_y:reset_n, settings_jerk_z:reset_n, settings_max_speed_e0:reset_n, settings_max_speed_e1:reset_n, settings_max_speed_x:reset_n, settings_max_speed_y:reset_n, settings_max_speed_z:reset_n, settings_max_temp_bed:reset_n, settings_max_temp_e0:reset_n, settings_max_temp_e1:reset_n, step_e0_now:reset_n, step_e1_now:reset_n, step_x_now:reset_n, step_y_now:reset_n, step_z_now:reset_n, sysid_qsys:reset_n, temp_0:reset_n, temp_1:reset_n, temp_2:reset_n, timing_e0_0:reset_n, timing_e0_1:reset_n, timing_e0_2:reset_n, timing_e0_3:reset_n, timing_e1_0:reset_n, timing_e1_1:reset_n, timing_e1_2:reset_n, timing_e1_3:reset_n, timing_x_0:reset_n, timing_x_1:reset_n, timing_x_2:reset_n, timing_x_3:reset_n, timing_y_0:reset_n, timing_y_1:reset_n, timing_y_2:reset_n, timing_y_3:reset_n, timing_z_0:reset_n, timing_z_1:reset_n, timing_z_2:reset_n, timing_z_3:reset_n]
	wire          rst_controller_001_reset_out_reset;                        // rst_controller_001:reset_out -> [mm_interconnect_0:hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_2:hps_0_f2h_axi_slave_agent_reset_sink_reset_bridge_in_reset_reset, mm_interconnect_3:hps_0_f2h_sdram0_data_translator_reset_reset_bridge_in_reset_reset]

	interrupt_latency_counter #(
		.INTR_TYPE    (0),
		.CLOCK_RATE   (50000000),
		.IRQ_PORT_CNT (3)
	) ilc (
		.reset_n     (~rst_controller_reset_out_reset),              //      reset_n.reset_n
		.clk         (clk_clk),                                      //          clk.clk
		.irq         (ilc_irq_irq),                                  //          irq.irq
		.avmm_addr   (mm_interconnect_1_ilc_avalon_slave_address),   // avalon_slave.address
		.avmm_wrdata (mm_interconnect_1_ilc_avalon_slave_writedata), //             .writedata
		.avmm_write  (mm_interconnect_1_ilc_avalon_slave_write),     //             .write
		.avmm_read   (mm_interconnect_1_ilc_avalon_slave_read),      //             .read
		.avmm_rddata (mm_interconnect_1_ilc_avalon_slave_readdata)   //             .readdata
	);

	soc_system_command_dt command_dt (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_1_command_dt_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_command_dt_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_command_dt_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_command_dt_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_command_dt_s1_readdata),   //                    .readdata
		.out_port   (command_dt_external_connection_export)       // external_connection.export
	);

	soc_system_command_e0 command_e0 (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_1_command_e0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_command_e0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_command_e0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_command_e0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_command_e0_s1_readdata),   //                    .readdata
		.out_port   (command_e0_external_connection_export)       // external_connection.export
	);

	soc_system_command_e0 command_e1 (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_1_command_e1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_command_e1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_command_e1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_command_e1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_command_e1_s1_readdata),   //                    .readdata
		.out_port   (command_e1_external_connection_export)       // external_connection.export
	);

	soc_system_command_e0 command_f_e0 (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_1_command_f_e0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_command_f_e0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_command_f_e0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_command_f_e0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_command_f_e0_s1_readdata),   //                    .readdata
		.out_port   (command_f_e0_external_connection_export)       // external_connection.export
	);

	soc_system_command_e0 command_f_e1 (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_1_command_f_e1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_command_f_e1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_command_f_e1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_command_f_e1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_command_f_e1_s1_readdata),   //                    .readdata
		.out_port   (command_f_e1_external_connection_export)       // external_connection.export
	);

	soc_system_command_e0 command_f_x (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_1_command_f_x_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_command_f_x_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_command_f_x_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_command_f_x_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_command_f_x_s1_readdata),   //                    .readdata
		.out_port   (command_f_x_external_connection_export)       // external_connection.export
	);

	soc_system_command_e0 command_f_y (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_1_command_f_y_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_command_f_y_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_command_f_y_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_command_f_y_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_command_f_y_s1_readdata),   //                    .readdata
		.out_port   (command_f_y_external_connection_export)       // external_connection.export
	);

	soc_system_command_e0 command_f_z (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_1_command_f_z_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_command_f_z_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_command_f_z_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_command_f_z_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_command_f_z_s1_readdata),   //                    .readdata
		.out_port   (command_f_z_external_connection_export)       // external_connection.export
	);

	soc_system_command_dt command_t (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_1_command_t_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_command_t_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_command_t_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_command_t_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_command_t_s1_readdata),   //                    .readdata
		.out_port   (command_t_external_connection_export)       // external_connection.export
	);

	soc_system_command_e0 command_type (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_1_command_type_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_command_type_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_command_type_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_command_type_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_command_type_s1_readdata),   //                    .readdata
		.out_port   (command_type_external_connection_export)       // external_connection.export
	);

	soc_system_command_e0 command_x (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_1_command_x_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_command_x_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_command_x_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_command_x_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_command_x_s1_readdata),   //                    .readdata
		.out_port   (command_x_external_connection_export)       // external_connection.export
	);

	soc_system_command_e0 command_y (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_1_command_y_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_command_y_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_command_y_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_command_y_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_command_y_s1_readdata),   //                    .readdata
		.out_port   (command_y_external_connection_export)       // external_connection.export
	);

	soc_system_command_e0 command_z (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_1_command_z_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_command_z_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_command_z_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_command_z_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_command_z_s1_readdata),   //                    .readdata
		.out_port   (command_z_external_connection_export)       // external_connection.export
	);

	soc_system_f2sdram_only_master #(
		.USE_PLI     (0),
		.PLI_PORT    (50000),
		.FIFO_DEPTHS (2)
	) f2sdram_only_master (
		.clk_clk              (clk_clk),                                  //          clk.clk
		.clk_reset_reset      (~reset_reset_n),                           //    clk_reset.reset
		.master_address       (f2sdram_only_master_master_address),       //       master.address
		.master_readdata      (f2sdram_only_master_master_readdata),      //             .readdata
		.master_read          (f2sdram_only_master_master_read),          //             .read
		.master_write         (f2sdram_only_master_master_write),         //             .write
		.master_writedata     (f2sdram_only_master_master_writedata),     //             .writedata
		.master_waitrequest   (f2sdram_only_master_master_waitrequest),   //             .waitrequest
		.master_readdatavalid (f2sdram_only_master_master_readdatavalid), //             .readdatavalid
		.master_byteenable    (f2sdram_only_master_master_byteenable),    //             .byteenable
		.master_reset_reset   ()                                          // master_reset.reset
	);

	soc_system_flags_in flags_in (
		.clk      (clk_clk),                                //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address  (mm_interconnect_1_flags_in_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_flags_in_s1_readdata), //                    .readdata
		.in_port  (flags_in_external_connection_export)     // external_connection.export
	);

	soc_system_command_e0 flags_out (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_1_flags_out_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_flags_out_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_flags_out_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_flags_out_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_flags_out_s1_readdata),   //                    .readdata
		.out_port   (flags_out_external_connection_export)       // external_connection.export
	);

	soc_system_f2sdram_only_master #(
		.USE_PLI     (0),
		.PLI_PORT    (50000),
		.FIFO_DEPTHS (2)
	) fpga_only_master (
		.clk_clk              (clk_clk),                               //          clk.clk
		.clk_reset_reset      (~reset_reset_n),                        //    clk_reset.reset
		.master_address       (fpga_only_master_master_address),       //       master.address
		.master_readdata      (fpga_only_master_master_readdata),      //             .readdata
		.master_read          (fpga_only_master_master_read),          //             .read
		.master_write         (fpga_only_master_master_write),         //             .write
		.master_writedata     (fpga_only_master_master_writedata),     //             .writedata
		.master_waitrequest   (fpga_only_master_master_waitrequest),   //             .waitrequest
		.master_readdatavalid (fpga_only_master_master_readdatavalid), //             .readdatavalid
		.master_byteenable    (fpga_only_master_master_byteenable),    //             .byteenable
		.master_reset_reset   ()                                       // master_reset.reset
	);

	soc_system_hps_0 #(
		.F2S_Width (2),
		.S2F_Width (2)
	) hps_0 (
		.f2h_cold_rst_req_n       (hps_0_f2h_cold_reset_req_reset_n),                      //  f2h_cold_reset_req.reset_n
		.f2h_dbg_rst_req_n        (hps_0_f2h_debug_reset_req_reset_n),                     // f2h_debug_reset_req.reset_n
		.f2h_warm_rst_req_n       (hps_0_f2h_warm_reset_req_reset_n),                      //  f2h_warm_reset_req.reset_n
		.f2h_stm_hwevents         (hps_0_f2h_stm_hw_events_stm_hwevents),                  //   f2h_stm_hw_events.stm_hwevents
		.uart1_cts                (hps_0_uart1_cts),                                       //               uart1.cts
		.uart1_dsr                (hps_0_uart1_dsr),                                       //                    .dsr
		.uart1_dcd                (hps_0_uart1_dcd),                                       //                    .dcd
		.uart1_ri                 (hps_0_uart1_ri),                                        //                    .ri
		.uart1_dtr                (hps_0_uart1_dtr),                                       //                    .dtr
		.uart1_rts                (hps_0_uart1_rts),                                       //                    .rts
		.uart1_out1_n             (hps_0_uart1_out1_n),                                    //                    .out1_n
		.uart1_out2_n             (hps_0_uart1_out2_n),                                    //                    .out2_n
		.uart1_rxd                (hps_0_uart1_rxd),                                       //                    .rxd
		.uart1_txd                (hps_0_uart1_txd),                                       //                    .txd
		.mem_a                    (memory_mem_a),                                          //              memory.mem_a
		.mem_ba                   (memory_mem_ba),                                         //                    .mem_ba
		.mem_ck                   (memory_mem_ck),                                         //                    .mem_ck
		.mem_ck_n                 (memory_mem_ck_n),                                       //                    .mem_ck_n
		.mem_cke                  (memory_mem_cke),                                        //                    .mem_cke
		.mem_cs_n                 (memory_mem_cs_n),                                       //                    .mem_cs_n
		.mem_ras_n                (memory_mem_ras_n),                                      //                    .mem_ras_n
		.mem_cas_n                (memory_mem_cas_n),                                      //                    .mem_cas_n
		.mem_we_n                 (memory_mem_we_n),                                       //                    .mem_we_n
		.mem_reset_n              (memory_mem_reset_n),                                    //                    .mem_reset_n
		.mem_dq                   (memory_mem_dq),                                         //                    .mem_dq
		.mem_dqs                  (memory_mem_dqs),                                        //                    .mem_dqs
		.mem_dqs_n                (memory_mem_dqs_n),                                      //                    .mem_dqs_n
		.mem_odt                  (memory_mem_odt),                                        //                    .mem_odt
		.mem_dm                   (memory_mem_dm),                                         //                    .mem_dm
		.oct_rzqin                (memory_oct_rzqin),                                      //                    .oct_rzqin
		.hps_io_emac1_inst_TX_CLK (hps_0_hps_io_hps_io_emac1_inst_TX_CLK),                 //              hps_io.hps_io_emac1_inst_TX_CLK
		.hps_io_emac1_inst_TXD0   (hps_0_hps_io_hps_io_emac1_inst_TXD0),                   //                    .hps_io_emac1_inst_TXD0
		.hps_io_emac1_inst_TXD1   (hps_0_hps_io_hps_io_emac1_inst_TXD1),                   //                    .hps_io_emac1_inst_TXD1
		.hps_io_emac1_inst_TXD2   (hps_0_hps_io_hps_io_emac1_inst_TXD2),                   //                    .hps_io_emac1_inst_TXD2
		.hps_io_emac1_inst_TXD3   (hps_0_hps_io_hps_io_emac1_inst_TXD3),                   //                    .hps_io_emac1_inst_TXD3
		.hps_io_emac1_inst_RXD0   (hps_0_hps_io_hps_io_emac1_inst_RXD0),                   //                    .hps_io_emac1_inst_RXD0
		.hps_io_emac1_inst_MDIO   (hps_0_hps_io_hps_io_emac1_inst_MDIO),                   //                    .hps_io_emac1_inst_MDIO
		.hps_io_emac1_inst_MDC    (hps_0_hps_io_hps_io_emac1_inst_MDC),                    //                    .hps_io_emac1_inst_MDC
		.hps_io_emac1_inst_RX_CTL (hps_0_hps_io_hps_io_emac1_inst_RX_CTL),                 //                    .hps_io_emac1_inst_RX_CTL
		.hps_io_emac1_inst_TX_CTL (hps_0_hps_io_hps_io_emac1_inst_TX_CTL),                 //                    .hps_io_emac1_inst_TX_CTL
		.hps_io_emac1_inst_RX_CLK (hps_0_hps_io_hps_io_emac1_inst_RX_CLK),                 //                    .hps_io_emac1_inst_RX_CLK
		.hps_io_emac1_inst_RXD1   (hps_0_hps_io_hps_io_emac1_inst_RXD1),                   //                    .hps_io_emac1_inst_RXD1
		.hps_io_emac1_inst_RXD2   (hps_0_hps_io_hps_io_emac1_inst_RXD2),                   //                    .hps_io_emac1_inst_RXD2
		.hps_io_emac1_inst_RXD3   (hps_0_hps_io_hps_io_emac1_inst_RXD3),                   //                    .hps_io_emac1_inst_RXD3
		.hps_io_sdio_inst_CMD     (hps_0_hps_io_hps_io_sdio_inst_CMD),                     //                    .hps_io_sdio_inst_CMD
		.hps_io_sdio_inst_D0      (hps_0_hps_io_hps_io_sdio_inst_D0),                      //                    .hps_io_sdio_inst_D0
		.hps_io_sdio_inst_D1      (hps_0_hps_io_hps_io_sdio_inst_D1),                      //                    .hps_io_sdio_inst_D1
		.hps_io_sdio_inst_CLK     (hps_0_hps_io_hps_io_sdio_inst_CLK),                     //                    .hps_io_sdio_inst_CLK
		.hps_io_sdio_inst_D2      (hps_0_hps_io_hps_io_sdio_inst_D2),                      //                    .hps_io_sdio_inst_D2
		.hps_io_sdio_inst_D3      (hps_0_hps_io_hps_io_sdio_inst_D3),                      //                    .hps_io_sdio_inst_D3
		.hps_io_usb1_inst_D0      (hps_0_hps_io_hps_io_usb1_inst_D0),                      //                    .hps_io_usb1_inst_D0
		.hps_io_usb1_inst_D1      (hps_0_hps_io_hps_io_usb1_inst_D1),                      //                    .hps_io_usb1_inst_D1
		.hps_io_usb1_inst_D2      (hps_0_hps_io_hps_io_usb1_inst_D2),                      //                    .hps_io_usb1_inst_D2
		.hps_io_usb1_inst_D3      (hps_0_hps_io_hps_io_usb1_inst_D3),                      //                    .hps_io_usb1_inst_D3
		.hps_io_usb1_inst_D4      (hps_0_hps_io_hps_io_usb1_inst_D4),                      //                    .hps_io_usb1_inst_D4
		.hps_io_usb1_inst_D5      (hps_0_hps_io_hps_io_usb1_inst_D5),                      //                    .hps_io_usb1_inst_D5
		.hps_io_usb1_inst_D6      (hps_0_hps_io_hps_io_usb1_inst_D6),                      //                    .hps_io_usb1_inst_D6
		.hps_io_usb1_inst_D7      (hps_0_hps_io_hps_io_usb1_inst_D7),                      //                    .hps_io_usb1_inst_D7
		.hps_io_usb1_inst_CLK     (hps_0_hps_io_hps_io_usb1_inst_CLK),                     //                    .hps_io_usb1_inst_CLK
		.hps_io_usb1_inst_STP     (hps_0_hps_io_hps_io_usb1_inst_STP),                     //                    .hps_io_usb1_inst_STP
		.hps_io_usb1_inst_DIR     (hps_0_hps_io_hps_io_usb1_inst_DIR),                     //                    .hps_io_usb1_inst_DIR
		.hps_io_usb1_inst_NXT     (hps_0_hps_io_hps_io_usb1_inst_NXT),                     //                    .hps_io_usb1_inst_NXT
		.hps_io_spim1_inst_CLK    (hps_0_hps_io_hps_io_spim1_inst_CLK),                    //                    .hps_io_spim1_inst_CLK
		.hps_io_spim1_inst_MOSI   (hps_0_hps_io_hps_io_spim1_inst_MOSI),                   //                    .hps_io_spim1_inst_MOSI
		.hps_io_spim1_inst_MISO   (hps_0_hps_io_hps_io_spim1_inst_MISO),                   //                    .hps_io_spim1_inst_MISO
		.hps_io_spim1_inst_SS0    (hps_0_hps_io_hps_io_spim1_inst_SS0),                    //                    .hps_io_spim1_inst_SS0
		.hps_io_uart0_inst_RX     (hps_0_hps_io_hps_io_uart0_inst_RX),                     //                    .hps_io_uart0_inst_RX
		.hps_io_uart0_inst_TX     (hps_0_hps_io_hps_io_uart0_inst_TX),                     //                    .hps_io_uart0_inst_TX
		.hps_io_i2c0_inst_SDA     (hps_0_hps_io_hps_io_i2c0_inst_SDA),                     //                    .hps_io_i2c0_inst_SDA
		.hps_io_i2c0_inst_SCL     (hps_0_hps_io_hps_io_i2c0_inst_SCL),                     //                    .hps_io_i2c0_inst_SCL
		.hps_io_i2c1_inst_SDA     (hps_0_hps_io_hps_io_i2c1_inst_SDA),                     //                    .hps_io_i2c1_inst_SDA
		.hps_io_i2c1_inst_SCL     (hps_0_hps_io_hps_io_i2c1_inst_SCL),                     //                    .hps_io_i2c1_inst_SCL
		.hps_io_gpio_inst_GPIO09  (hps_0_hps_io_hps_io_gpio_inst_GPIO09),                  //                    .hps_io_gpio_inst_GPIO09
		.hps_io_gpio_inst_GPIO35  (hps_0_hps_io_hps_io_gpio_inst_GPIO35),                  //                    .hps_io_gpio_inst_GPIO35
		.hps_io_gpio_inst_GPIO40  (hps_0_hps_io_hps_io_gpio_inst_GPIO40),                  //                    .hps_io_gpio_inst_GPIO40
		.hps_io_gpio_inst_GPIO53  (hps_0_hps_io_hps_io_gpio_inst_GPIO53),                  //                    .hps_io_gpio_inst_GPIO53
		.hps_io_gpio_inst_GPIO54  (hps_0_hps_io_hps_io_gpio_inst_GPIO54),                  //                    .hps_io_gpio_inst_GPIO54
		.hps_io_gpio_inst_GPIO61  (hps_0_hps_io_hps_io_gpio_inst_GPIO61),                  //                    .hps_io_gpio_inst_GPIO61
		.h2f_rst_n                (hps_0_h2f_reset_reset_n),                               //           h2f_reset.reset_n
		.f2h_sdram0_clk           (clk_clk),                                               //    f2h_sdram0_clock.clk
		.f2h_sdram0_ADDRESS       (mm_interconnect_3_hps_0_f2h_sdram0_data_address),       //     f2h_sdram0_data.address
		.f2h_sdram0_BURSTCOUNT    (mm_interconnect_3_hps_0_f2h_sdram0_data_burstcount),    //                    .burstcount
		.f2h_sdram0_WAITREQUEST   (mm_interconnect_3_hps_0_f2h_sdram0_data_waitrequest),   //                    .waitrequest
		.f2h_sdram0_READDATA      (mm_interconnect_3_hps_0_f2h_sdram0_data_readdata),      //                    .readdata
		.f2h_sdram0_READDATAVALID (mm_interconnect_3_hps_0_f2h_sdram0_data_readdatavalid), //                    .readdatavalid
		.f2h_sdram0_READ          (mm_interconnect_3_hps_0_f2h_sdram0_data_read),          //                    .read
		.f2h_sdram0_WRITEDATA     (mm_interconnect_3_hps_0_f2h_sdram0_data_writedata),     //                    .writedata
		.f2h_sdram0_BYTEENABLE    (mm_interconnect_3_hps_0_f2h_sdram0_data_byteenable),    //                    .byteenable
		.f2h_sdram0_WRITE         (mm_interconnect_3_hps_0_f2h_sdram0_data_write),         //                    .write
		.h2f_axi_clk              (clk_clk),                                               //       h2f_axi_clock.clk
		.h2f_AWID                 (),                                                      //      h2f_axi_master.awid
		.h2f_AWADDR               (),                                                      //                    .awaddr
		.h2f_AWLEN                (),                                                      //                    .awlen
		.h2f_AWSIZE               (),                                                      //                    .awsize
		.h2f_AWBURST              (),                                                      //                    .awburst
		.h2f_AWLOCK               (),                                                      //                    .awlock
		.h2f_AWCACHE              (),                                                      //                    .awcache
		.h2f_AWPROT               (),                                                      //                    .awprot
		.h2f_AWVALID              (),                                                      //                    .awvalid
		.h2f_AWREADY              (),                                                      //                    .awready
		.h2f_WID                  (),                                                      //                    .wid
		.h2f_WDATA                (),                                                      //                    .wdata
		.h2f_WSTRB                (),                                                      //                    .wstrb
		.h2f_WLAST                (),                                                      //                    .wlast
		.h2f_WVALID               (),                                                      //                    .wvalid
		.h2f_WREADY               (),                                                      //                    .wready
		.h2f_BID                  (),                                                      //                    .bid
		.h2f_BRESP                (),                                                      //                    .bresp
		.h2f_BVALID               (),                                                      //                    .bvalid
		.h2f_BREADY               (),                                                      //                    .bready
		.h2f_ARID                 (),                                                      //                    .arid
		.h2f_ARADDR               (),                                                      //                    .araddr
		.h2f_ARLEN                (),                                                      //                    .arlen
		.h2f_ARSIZE               (),                                                      //                    .arsize
		.h2f_ARBURST              (),                                                      //                    .arburst
		.h2f_ARLOCK               (),                                                      //                    .arlock
		.h2f_ARCACHE              (),                                                      //                    .arcache
		.h2f_ARPROT               (),                                                      //                    .arprot
		.h2f_ARVALID              (),                                                      //                    .arvalid
		.h2f_ARREADY              (),                                                      //                    .arready
		.h2f_RID                  (),                                                      //                    .rid
		.h2f_RDATA                (),                                                      //                    .rdata
		.h2f_RRESP                (),                                                      //                    .rresp
		.h2f_RLAST                (),                                                      //                    .rlast
		.h2f_RVALID               (),                                                      //                    .rvalid
		.h2f_RREADY               (),                                                      //                    .rready
		.f2h_axi_clk              (clk_clk),                                               //       f2h_axi_clock.clk
		.f2h_AWID                 (mm_interconnect_2_hps_0_f2h_axi_slave_awid),            //       f2h_axi_slave.awid
		.f2h_AWADDR               (mm_interconnect_2_hps_0_f2h_axi_slave_awaddr),          //                    .awaddr
		.f2h_AWLEN                (mm_interconnect_2_hps_0_f2h_axi_slave_awlen),           //                    .awlen
		.f2h_AWSIZE               (mm_interconnect_2_hps_0_f2h_axi_slave_awsize),          //                    .awsize
		.f2h_AWBURST              (mm_interconnect_2_hps_0_f2h_axi_slave_awburst),         //                    .awburst
		.f2h_AWLOCK               (mm_interconnect_2_hps_0_f2h_axi_slave_awlock),          //                    .awlock
		.f2h_AWCACHE              (mm_interconnect_2_hps_0_f2h_axi_slave_awcache),         //                    .awcache
		.f2h_AWPROT               (mm_interconnect_2_hps_0_f2h_axi_slave_awprot),          //                    .awprot
		.f2h_AWVALID              (mm_interconnect_2_hps_0_f2h_axi_slave_awvalid),         //                    .awvalid
		.f2h_AWREADY              (mm_interconnect_2_hps_0_f2h_axi_slave_awready),         //                    .awready
		.f2h_AWUSER               (mm_interconnect_2_hps_0_f2h_axi_slave_awuser),          //                    .awuser
		.f2h_WID                  (mm_interconnect_2_hps_0_f2h_axi_slave_wid),             //                    .wid
		.f2h_WDATA                (mm_interconnect_2_hps_0_f2h_axi_slave_wdata),           //                    .wdata
		.f2h_WSTRB                (mm_interconnect_2_hps_0_f2h_axi_slave_wstrb),           //                    .wstrb
		.f2h_WLAST                (mm_interconnect_2_hps_0_f2h_axi_slave_wlast),           //                    .wlast
		.f2h_WVALID               (mm_interconnect_2_hps_0_f2h_axi_slave_wvalid),          //                    .wvalid
		.f2h_WREADY               (mm_interconnect_2_hps_0_f2h_axi_slave_wready),          //                    .wready
		.f2h_BID                  (mm_interconnect_2_hps_0_f2h_axi_slave_bid),             //                    .bid
		.f2h_BRESP                (mm_interconnect_2_hps_0_f2h_axi_slave_bresp),           //                    .bresp
		.f2h_BVALID               (mm_interconnect_2_hps_0_f2h_axi_slave_bvalid),          //                    .bvalid
		.f2h_BREADY               (mm_interconnect_2_hps_0_f2h_axi_slave_bready),          //                    .bready
		.f2h_ARID                 (mm_interconnect_2_hps_0_f2h_axi_slave_arid),            //                    .arid
		.f2h_ARADDR               (mm_interconnect_2_hps_0_f2h_axi_slave_araddr),          //                    .araddr
		.f2h_ARLEN                (mm_interconnect_2_hps_0_f2h_axi_slave_arlen),           //                    .arlen
		.f2h_ARSIZE               (mm_interconnect_2_hps_0_f2h_axi_slave_arsize),          //                    .arsize
		.f2h_ARBURST              (mm_interconnect_2_hps_0_f2h_axi_slave_arburst),         //                    .arburst
		.f2h_ARLOCK               (mm_interconnect_2_hps_0_f2h_axi_slave_arlock),          //                    .arlock
		.f2h_ARCACHE              (mm_interconnect_2_hps_0_f2h_axi_slave_arcache),         //                    .arcache
		.f2h_ARPROT               (mm_interconnect_2_hps_0_f2h_axi_slave_arprot),          //                    .arprot
		.f2h_ARVALID              (mm_interconnect_2_hps_0_f2h_axi_slave_arvalid),         //                    .arvalid
		.f2h_ARREADY              (mm_interconnect_2_hps_0_f2h_axi_slave_arready),         //                    .arready
		.f2h_ARUSER               (mm_interconnect_2_hps_0_f2h_axi_slave_aruser),          //                    .aruser
		.f2h_RID                  (mm_interconnect_2_hps_0_f2h_axi_slave_rid),             //                    .rid
		.f2h_RDATA                (mm_interconnect_2_hps_0_f2h_axi_slave_rdata),           //                    .rdata
		.f2h_RRESP                (mm_interconnect_2_hps_0_f2h_axi_slave_rresp),           //                    .rresp
		.f2h_RLAST                (mm_interconnect_2_hps_0_f2h_axi_slave_rlast),           //                    .rlast
		.f2h_RVALID               (mm_interconnect_2_hps_0_f2h_axi_slave_rvalid),          //                    .rvalid
		.f2h_RREADY               (mm_interconnect_2_hps_0_f2h_axi_slave_rready),          //                    .rready
		.h2f_lw_axi_clk           (clk_clk),                                               //    h2f_lw_axi_clock.clk
		.h2f_lw_AWID              (hps_0_h2f_lw_axi_master_awid),                          //   h2f_lw_axi_master.awid
		.h2f_lw_AWADDR            (hps_0_h2f_lw_axi_master_awaddr),                        //                    .awaddr
		.h2f_lw_AWLEN             (hps_0_h2f_lw_axi_master_awlen),                         //                    .awlen
		.h2f_lw_AWSIZE            (hps_0_h2f_lw_axi_master_awsize),                        //                    .awsize
		.h2f_lw_AWBURST           (hps_0_h2f_lw_axi_master_awburst),                       //                    .awburst
		.h2f_lw_AWLOCK            (hps_0_h2f_lw_axi_master_awlock),                        //                    .awlock
		.h2f_lw_AWCACHE           (hps_0_h2f_lw_axi_master_awcache),                       //                    .awcache
		.h2f_lw_AWPROT            (hps_0_h2f_lw_axi_master_awprot),                        //                    .awprot
		.h2f_lw_AWVALID           (hps_0_h2f_lw_axi_master_awvalid),                       //                    .awvalid
		.h2f_lw_AWREADY           (hps_0_h2f_lw_axi_master_awready),                       //                    .awready
		.h2f_lw_WID               (hps_0_h2f_lw_axi_master_wid),                           //                    .wid
		.h2f_lw_WDATA             (hps_0_h2f_lw_axi_master_wdata),                         //                    .wdata
		.h2f_lw_WSTRB             (hps_0_h2f_lw_axi_master_wstrb),                         //                    .wstrb
		.h2f_lw_WLAST             (hps_0_h2f_lw_axi_master_wlast),                         //                    .wlast
		.h2f_lw_WVALID            (hps_0_h2f_lw_axi_master_wvalid),                        //                    .wvalid
		.h2f_lw_WREADY            (hps_0_h2f_lw_axi_master_wready),                        //                    .wready
		.h2f_lw_BID               (hps_0_h2f_lw_axi_master_bid),                           //                    .bid
		.h2f_lw_BRESP             (hps_0_h2f_lw_axi_master_bresp),                         //                    .bresp
		.h2f_lw_BVALID            (hps_0_h2f_lw_axi_master_bvalid),                        //                    .bvalid
		.h2f_lw_BREADY            (hps_0_h2f_lw_axi_master_bready),                        //                    .bready
		.h2f_lw_ARID              (hps_0_h2f_lw_axi_master_arid),                          //                    .arid
		.h2f_lw_ARADDR            (hps_0_h2f_lw_axi_master_araddr),                        //                    .araddr
		.h2f_lw_ARLEN             (hps_0_h2f_lw_axi_master_arlen),                         //                    .arlen
		.h2f_lw_ARSIZE            (hps_0_h2f_lw_axi_master_arsize),                        //                    .arsize
		.h2f_lw_ARBURST           (hps_0_h2f_lw_axi_master_arburst),                       //                    .arburst
		.h2f_lw_ARLOCK            (hps_0_h2f_lw_axi_master_arlock),                        //                    .arlock
		.h2f_lw_ARCACHE           (hps_0_h2f_lw_axi_master_arcache),                       //                    .arcache
		.h2f_lw_ARPROT            (hps_0_h2f_lw_axi_master_arprot),                        //                    .arprot
		.h2f_lw_ARVALID           (hps_0_h2f_lw_axi_master_arvalid),                       //                    .arvalid
		.h2f_lw_ARREADY           (hps_0_h2f_lw_axi_master_arready),                       //                    .arready
		.h2f_lw_RID               (hps_0_h2f_lw_axi_master_rid),                           //                    .rid
		.h2f_lw_RDATA             (hps_0_h2f_lw_axi_master_rdata),                         //                    .rdata
		.h2f_lw_RRESP             (hps_0_h2f_lw_axi_master_rresp),                         //                    .rresp
		.h2f_lw_RLAST             (hps_0_h2f_lw_axi_master_rlast),                         //                    .rlast
		.h2f_lw_RVALID            (hps_0_h2f_lw_axi_master_rvalid),                        //                    .rvalid
		.h2f_lw_RREADY            (hps_0_h2f_lw_axi_master_rready),                        //                    .rready
		.f2h_irq_p0               (hps_0_f2h_irq0_irq),                                    //            f2h_irq0.irq
		.f2h_irq_p1               (hps_0_f2h_irq1_irq)                                     //            f2h_irq1.irq
	);

	soc_system_f2sdram_only_master #(
		.USE_PLI     (0),
		.PLI_PORT    (50000),
		.FIFO_DEPTHS (2)
	) hps_only_master (
		.clk_clk              (clk_clk),                              //          clk.clk
		.clk_reset_reset      (~reset_reset_n),                       //    clk_reset.reset
		.master_address       (hps_only_master_master_address),       //       master.address
		.master_readdata      (hps_only_master_master_readdata),      //             .readdata
		.master_read          (hps_only_master_master_read),          //             .read
		.master_write         (hps_only_master_master_write),         //             .write
		.master_writedata     (hps_only_master_master_writedata),     //             .writedata
		.master_waitrequest   (hps_only_master_master_waitrequest),   //             .waitrequest
		.master_readdatavalid (hps_only_master_master_readdatavalid), //             .readdatavalid
		.master_byteenable    (hps_only_master_master_byteenable),    //             .byteenable
		.master_reset_reset   ()                                      // master_reset.reset
	);

	soc_system_jtag_uart jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_1_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_1_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_1_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                   //               irq.irq
	);

	soc_system_flags_in max_params_0 (
		.clk      (clk_clk),                                    //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address  (mm_interconnect_1_max_params_0_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_max_params_0_s1_readdata), //                    .readdata
		.in_port  (max_params_0_external_connection_export)     // external_connection.export
	);

	soc_system_flags_in max_params_1 (
		.clk      (clk_clk),                                    //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address  (mm_interconnect_1_max_params_1_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_max_params_1_s1_readdata), //                    .readdata
		.in_port  (max_params_1_external_connection_export)     // external_connection.export
	);

	soc_system_flags_in max_params_2 (
		.clk      (clk_clk),                                    //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address  (mm_interconnect_1_max_params_2_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_max_params_2_s1_readdata), //                    .readdata
		.in_port  (max_params_2_external_connection_export)     // external_connection.export
	);

	soc_system_flags_in max_params_3 (
		.clk      (clk_clk),                                    //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address  (mm_interconnect_1_max_params_3_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_max_params_3_s1_readdata), //                    .readdata
		.in_port  (max_params_3_external_connection_export)     // external_connection.export
	);

	soc_system_flags_in max_params_4 (
		.clk      (clk_clk),                                    //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address  (mm_interconnect_1_max_params_4_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_max_params_4_s1_readdata), //                    .readdata
		.in_port  (max_params_4_external_connection_export)     // external_connection.export
	);

	soc_system_flags_in max_timing_0 (
		.clk      (clk_clk),                                    //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address  (mm_interconnect_1_max_timing_0_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_max_timing_0_s1_readdata), //                    .readdata
		.in_port  (max_timing_0_external_connection_export)     // external_connection.export
	);

	soc_system_flags_in max_timing_1 (
		.clk      (clk_clk),                                    //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address  (mm_interconnect_1_max_timing_1_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_max_timing_1_s1_readdata), //                    .readdata
		.in_port  (max_timing_1_external_connection_export)     // external_connection.export
	);

	soc_system_flags_in max_timing_2 (
		.clk      (clk_clk),                                    //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address  (mm_interconnect_1_max_timing_2_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_max_timing_2_s1_readdata), //                    .readdata
		.in_port  (max_timing_2_external_connection_export)     // external_connection.export
	);

	soc_system_flags_in max_timing_3 (
		.clk      (clk_clk),                                    //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address  (mm_interconnect_1_max_timing_3_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_max_timing_3_s1_readdata), //                    .readdata
		.in_port  (max_timing_3_external_connection_export)     // external_connection.export
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (32),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (18),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) mm_bridge_0 (
		.clk              (clk_clk),                                        //   clk.clk
		.reset            (rst_controller_reset_out_reset),                 // reset.reset
		.s0_waitrequest   (mm_interconnect_0_mm_bridge_0_s0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (mm_interconnect_0_mm_bridge_0_s0_readdata),      //      .readdata
		.s0_readdatavalid (mm_interconnect_0_mm_bridge_0_s0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (mm_interconnect_0_mm_bridge_0_s0_burstcount),    //      .burstcount
		.s0_writedata     (mm_interconnect_0_mm_bridge_0_s0_writedata),     //      .writedata
		.s0_address       (mm_interconnect_0_mm_bridge_0_s0_address),       //      .address
		.s0_write         (mm_interconnect_0_mm_bridge_0_s0_write),         //      .write
		.s0_read          (mm_interconnect_0_mm_bridge_0_s0_read),          //      .read
		.s0_byteenable    (mm_interconnect_0_mm_bridge_0_s0_byteenable),    //      .byteenable
		.s0_debugaccess   (mm_interconnect_0_mm_bridge_0_s0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (mm_bridge_0_m0_waitrequest),                     //    m0.waitrequest
		.m0_readdata      (mm_bridge_0_m0_readdata),                        //      .readdata
		.m0_readdatavalid (mm_bridge_0_m0_readdatavalid),                   //      .readdatavalid
		.m0_burstcount    (mm_bridge_0_m0_burstcount),                      //      .burstcount
		.m0_writedata     (mm_bridge_0_m0_writedata),                       //      .writedata
		.m0_address       (mm_bridge_0_m0_address),                         //      .address
		.m0_write         (mm_bridge_0_m0_write),                           //      .write
		.m0_read          (mm_bridge_0_m0_read),                            //      .read
		.m0_byteenable    (mm_bridge_0_m0_byteenable),                      //      .byteenable
		.m0_debugaccess   (mm_bridge_0_m0_debugaccess),                     //      .debugaccess
		.s0_response      (),                                               // (terminated)
		.m0_response      (2'b00)                                           // (terminated)
	);

	soc_system_flags_in new_rparams_e0_0 (
		.clk      (clk_clk),                                        //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address  (mm_interconnect_1_new_rparams_e0_0_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_new_rparams_e0_0_s1_readdata), //                    .readdata
		.in_port  (new_rparams_e0_0_external_connection_export)     // external_connection.export
	);

	soc_system_flags_in new_rparams_e0_1 (
		.clk      (clk_clk),                                        //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address  (mm_interconnect_1_new_rparams_e0_1_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_new_rparams_e0_1_s1_readdata), //                    .readdata
		.in_port  (new_rparams_e0_1_external_connection_export)     // external_connection.export
	);

	soc_system_flags_in new_rparams_e0_2 (
		.clk      (clk_clk),                                        //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address  (mm_interconnect_1_new_rparams_e0_2_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_new_rparams_e0_2_s1_readdata), //                    .readdata
		.in_port  (new_rparams_e0_2_external_connection_export)     // external_connection.export
	);

	soc_system_flags_in new_rparams_e0_3 (
		.clk      (clk_clk),                                        //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address  (mm_interconnect_1_new_rparams_e0_3_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_new_rparams_e0_3_s1_readdata), //                    .readdata
		.in_port  (new_rparams_e0_3_external_connection_export)     // external_connection.export
	);

	soc_system_flags_in new_rparams_e0_4 (
		.clk      (clk_clk),                                        //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address  (mm_interconnect_1_new_rparams_e0_4_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_new_rparams_e0_4_s1_readdata), //                    .readdata
		.in_port  (new_rparams_e0_4_external_connection_export)     // external_connection.export
	);

	soc_system_flags_in new_rparams_e1_0 (
		.clk      (clk_clk),                                        //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address  (mm_interconnect_1_new_rparams_e1_0_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_new_rparams_e1_0_s1_readdata), //                    .readdata
		.in_port  (new_rparams_e1_0_external_connection_export)     // external_connection.export
	);

	soc_system_flags_in new_rparams_e1_1 (
		.clk      (clk_clk),                                        //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address  (mm_interconnect_1_new_rparams_e1_1_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_new_rparams_e1_1_s1_readdata), //                    .readdata
		.in_port  (new_rparams_e1_1_external_connection_export)     // external_connection.export
	);

	soc_system_flags_in new_rparams_e1_2 (
		.clk      (clk_clk),                                        //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address  (mm_interconnect_1_new_rparams_e1_2_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_new_rparams_e1_2_s1_readdata), //                    .readdata
		.in_port  (new_rparams_e1_2_external_connection_export)     // external_connection.export
	);

	soc_system_flags_in new_rparams_e1_3 (
		.clk      (clk_clk),                                        //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address  (mm_interconnect_1_new_rparams_e1_3_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_new_rparams_e1_3_s1_readdata), //                    .readdata
		.in_port  (new_rparams_e1_3_external_connection_export)     // external_connection.export
	);

	soc_system_flags_in new_rparams_e1_4 (
		.clk      (clk_clk),                                        //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address  (mm_interconnect_1_new_rparams_e1_4_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_new_rparams_e1_4_s1_readdata), //                    .readdata
		.in_port  (new_rparams_e1_4_external_connection_export)     // external_connection.export
	);

	soc_system_flags_in new_rparams_x_0 (
		.clk      (clk_clk),                                       //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address  (mm_interconnect_1_new_rparams_x_0_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_new_rparams_x_0_s1_readdata), //                    .readdata
		.in_port  (new_rparams_x_0_external_connection_export)     // external_connection.export
	);

	soc_system_flags_in new_rparams_x_1 (
		.clk      (clk_clk),                                       //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address  (mm_interconnect_1_new_rparams_x_1_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_new_rparams_x_1_s1_readdata), //                    .readdata
		.in_port  (new_rparams_x_1_external_connection_export)     // external_connection.export
	);

	soc_system_flags_in new_rparams_x_2 (
		.clk      (clk_clk),                                       //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address  (mm_interconnect_1_new_rparams_x_2_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_new_rparams_x_2_s1_readdata), //                    .readdata
		.in_port  (new_rparams_x_2_external_connection_export)     // external_connection.export
	);

	soc_system_flags_in new_rparams_x_3 (
		.clk      (clk_clk),                                       //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address  (mm_interconnect_1_new_rparams_x_3_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_new_rparams_x_3_s1_readdata), //                    .readdata
		.in_port  (new_rparams_x_3_external_connection_export)     // external_connection.export
	);

	soc_system_flags_in new_rparams_x_4 (
		.clk      (clk_clk),                                       //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address  (mm_interconnect_1_new_rparams_x_4_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_new_rparams_x_4_s1_readdata), //                    .readdata
		.in_port  (new_rparams_x_4_external_connection_export)     // external_connection.export
	);

	soc_system_flags_in new_rparams_y_0 (
		.clk      (clk_clk),                                       //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address  (mm_interconnect_1_new_rparams_y_0_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_new_rparams_y_0_s1_readdata), //                    .readdata
		.in_port  (new_rparams_y_0_external_connection_export)     // external_connection.export
	);

	soc_system_flags_in new_rparams_y_1 (
		.clk      (clk_clk),                                       //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address  (mm_interconnect_1_new_rparams_y_1_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_new_rparams_y_1_s1_readdata), //                    .readdata
		.in_port  (new_rparams_y_1_external_connection_export)     // external_connection.export
	);

	soc_system_flags_in new_rparams_y_2 (
		.clk      (clk_clk),                                       //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address  (mm_interconnect_1_new_rparams_y_2_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_new_rparams_y_2_s1_readdata), //                    .readdata
		.in_port  (new_rparams_y_2_external_connection_export)     // external_connection.export
	);

	soc_system_flags_in new_rparams_y_3 (
		.clk      (clk_clk),                                       //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address  (mm_interconnect_1_new_rparams_y_3_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_new_rparams_y_3_s1_readdata), //                    .readdata
		.in_port  (new_rparams_y_3_external_connection_export)     // external_connection.export
	);

	soc_system_flags_in new_rparams_y_4 (
		.clk      (clk_clk),                                       //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address  (mm_interconnect_1_new_rparams_y_4_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_new_rparams_y_4_s1_readdata), //                    .readdata
		.in_port  (new_rparams_y_4_external_connection_export)     // external_connection.export
	);

	soc_system_flags_in new_rparams_z_0 (
		.clk      (clk_clk),                                       //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address  (mm_interconnect_1_new_rparams_z_0_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_new_rparams_z_0_s1_readdata), //                    .readdata
		.in_port  (new_rparams_z_0_external_connection_export)     // external_connection.export
	);

	soc_system_flags_in new_rparams_z_1 (
		.clk      (clk_clk),                                       //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address  (mm_interconnect_1_new_rparams_z_1_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_new_rparams_z_1_s1_readdata), //                    .readdata
		.in_port  (new_rparams_z_1_external_connection_export)     // external_connection.export
	);

	soc_system_flags_in new_rparams_z_2 (
		.clk      (clk_clk),                                       //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address  (mm_interconnect_1_new_rparams_z_2_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_new_rparams_z_2_s1_readdata), //                    .readdata
		.in_port  (new_rparams_z_2_external_connection_export)     // external_connection.export
	);

	soc_system_flags_in new_rparams_z_3 (
		.clk      (clk_clk),                                       //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address  (mm_interconnect_1_new_rparams_z_3_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_new_rparams_z_3_s1_readdata), //                    .readdata
		.in_port  (new_rparams_z_3_external_connection_export)     // external_connection.export
	);

	soc_system_flags_in new_rparams_z_4 (
		.clk      (clk_clk),                                       //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address  (mm_interconnect_1_new_rparams_z_4_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_new_rparams_z_4_s1_readdata), //                    .readdata
		.in_port  (new_rparams_z_4_external_connection_export)     // external_connection.export
	);

	soc_system_flags_in params_e0_0 (
		.clk      (clk_clk),                                   //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address  (mm_interconnect_1_params_e0_0_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_params_e0_0_s1_readdata), //                    .readdata
		.in_port  (params_e0_0_external_connection_export)     // external_connection.export
	);

	soc_system_flags_in params_e0_1 (
		.clk      (clk_clk),                                   //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address  (mm_interconnect_1_params_e0_1_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_params_e0_1_s1_readdata), //                    .readdata
		.in_port  (params_e0_1_external_connection_export)     // external_connection.export
	);

	soc_system_flags_in params_e0_2 (
		.clk      (clk_clk),                                   //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address  (mm_interconnect_1_params_e0_2_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_params_e0_2_s1_readdata), //                    .readdata
		.in_port  (params_e0_2_external_connection_export)     // external_connection.export
	);

	soc_system_flags_in params_e0_3 (
		.clk      (clk_clk),                                   //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address  (mm_interconnect_1_params_e0_3_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_params_e0_3_s1_readdata), //                    .readdata
		.in_port  (params_e0_3_external_connection_export)     // external_connection.export
	);

	soc_system_flags_in params_e0_4 (
		.clk      (clk_clk),                                   //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address  (mm_interconnect_1_params_e0_4_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_params_e0_4_s1_readdata), //                    .readdata
		.in_port  (params_e0_4_external_connection_export)     // external_connection.export
	);

	soc_system_flags_in params_e1_0 (
		.clk      (clk_clk),                                   //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address  (mm_interconnect_1_params_e1_0_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_params_e1_0_s1_readdata), //                    .readdata
		.in_port  (params_e1_0_external_connection_export)     // external_connection.export
	);

	soc_system_flags_in params_e1_1 (
		.clk      (clk_clk),                                   //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address  (mm_interconnect_1_params_e1_1_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_params_e1_1_s1_readdata), //                    .readdata
		.in_port  (params_e1_1_external_connection_export)     // external_connection.export
	);

	soc_system_flags_in params_e1_2 (
		.clk      (clk_clk),                                   //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address  (mm_interconnect_1_params_e1_2_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_params_e1_2_s1_readdata), //                    .readdata
		.in_port  (params_e1_2_external_connection_export)     // external_connection.export
	);

	soc_system_flags_in params_e1_3 (
		.clk      (clk_clk),                                   //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address  (mm_interconnect_1_params_e1_3_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_params_e1_3_s1_readdata), //                    .readdata
		.in_port  (params_e1_3_external_connection_export)     // external_connection.export
	);

	soc_system_flags_in params_e1_4 (
		.clk      (clk_clk),                                   //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address  (mm_interconnect_1_params_e1_4_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_params_e1_4_s1_readdata), //                    .readdata
		.in_port  (params_e1_4_external_connection_export)     // external_connection.export
	);

	soc_system_flags_in params_x_0 (
		.clk      (clk_clk),                                  //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_1_params_x_0_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_params_x_0_s1_readdata), //                    .readdata
		.in_port  (params_x_0_external_connection_export)     // external_connection.export
	);

	soc_system_flags_in params_x_1 (
		.clk      (clk_clk),                                  //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_1_params_x_1_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_params_x_1_s1_readdata), //                    .readdata
		.in_port  (params_x_1_external_connection_export)     // external_connection.export
	);

	soc_system_flags_in params_x_2 (
		.clk      (clk_clk),                                  //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_1_params_x_2_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_params_x_2_s1_readdata), //                    .readdata
		.in_port  (params_x_2_external_connection_export)     // external_connection.export
	);

	soc_system_flags_in params_x_3 (
		.clk      (clk_clk),                                  //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_1_params_x_3_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_params_x_3_s1_readdata), //                    .readdata
		.in_port  (params_x_3_external_connection_export)     // external_connection.export
	);

	soc_system_flags_in params_x_4 (
		.clk      (clk_clk),                                  //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_1_params_x_4_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_params_x_4_s1_readdata), //                    .readdata
		.in_port  (params_x_4_external_connection_export)     // external_connection.export
	);

	soc_system_flags_in params_y_0 (
		.clk      (clk_clk),                                  //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_1_params_y_0_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_params_y_0_s1_readdata), //                    .readdata
		.in_port  (params_y_0_external_connection_export)     // external_connection.export
	);

	soc_system_flags_in params_y_1 (
		.clk      (clk_clk),                                  //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_1_params_y_1_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_params_y_1_s1_readdata), //                    .readdata
		.in_port  (params_y_1_external_connection_export)     // external_connection.export
	);

	soc_system_flags_in params_y_2 (
		.clk      (clk_clk),                                  //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_1_params_y_2_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_params_y_2_s1_readdata), //                    .readdata
		.in_port  (params_y_2_external_connection_export)     // external_connection.export
	);

	soc_system_flags_in params_y_3 (
		.clk      (clk_clk),                                  //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_1_params_y_3_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_params_y_3_s1_readdata), //                    .readdata
		.in_port  (params_y_3_external_connection_export)     // external_connection.export
	);

	soc_system_flags_in params_y_4 (
		.clk      (clk_clk),                                  //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_1_params_y_4_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_params_y_4_s1_readdata), //                    .readdata
		.in_port  (params_y_4_external_connection_export)     // external_connection.export
	);

	soc_system_flags_in params_z_0 (
		.clk      (clk_clk),                                  //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_1_params_z_0_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_params_z_0_s1_readdata), //                    .readdata
		.in_port  (params_z_0_external_connection_export)     // external_connection.export
	);

	soc_system_flags_in params_z_1 (
		.clk      (clk_clk),                                  //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_1_params_z_1_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_params_z_1_s1_readdata), //                    .readdata
		.in_port  (params_z_1_external_connection_export)     // external_connection.export
	);

	soc_system_flags_in params_z_2 (
		.clk      (clk_clk),                                  //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_1_params_z_2_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_params_z_2_s1_readdata), //                    .readdata
		.in_port  (params_z_2_external_connection_export)     // external_connection.export
	);

	soc_system_flags_in params_z_3 (
		.clk      (clk_clk),                                  //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_1_params_z_3_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_params_z_3_s1_readdata), //                    .readdata
		.in_port  (params_z_3_external_connection_export)     // external_connection.export
	);

	soc_system_flags_in params_z_4 (
		.clk      (clk_clk),                                  //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_1_params_z_4_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_params_z_4_s1_readdata), //                    .readdata
		.in_port  (params_z_4_external_connection_export)     // external_connection.export
	);

	soc_system_pll_sys pll_sys (
		.refclk   (clk_clk),                  //  refclk.clk
		.rst      (~reset_reset_n),           //   reset.reset
		.outclk_0 (pll_sys_outclk100mhz_clk), // outclk0.clk
		.outclk_1 (pll_sys_outclk10mhz_clk),  // outclk1.clk
		.outclk_2 (pll_sys_outclk5mhz_clk),   // outclk2.clk
		.outclk_3 (pll_sys_outclk1mhz_clk),   // outclk3.clk
		.locked   ()                          // (terminated)
	);

	soc_system_position_e0 position_e0 (
		.clk      (clk_clk),                                   //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address  (mm_interconnect_1_position_e0_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_position_e0_s1_readdata), //                    .readdata
		.in_port  (position_e0_external_connection_export)     // external_connection.export
	);

	soc_system_position_e0 position_e1 (
		.clk      (clk_clk),                                   //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address  (mm_interconnect_1_position_e1_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_position_e1_s1_readdata), //                    .readdata
		.in_port  (position_e1_external_connection_export)     // external_connection.export
	);

	soc_system_position_e0 position_x (
		.clk      (clk_clk),                                  //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_1_position_x_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_position_x_s1_readdata), //                    .readdata
		.in_port  (position_x_external_connection_export)     // external_connection.export
	);

	soc_system_position_e0 position_y (
		.clk      (clk_clk),                                  //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_1_position_y_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_position_y_s1_readdata), //                    .readdata
		.in_port  (position_y_external_connection_export)     // external_connection.export
	);

	soc_system_position_e0 position_z (
		.clk      (clk_clk),                                  //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_1_position_z_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_position_z_s1_readdata), //                    .readdata
		.in_port  (position_z_external_connection_export)     // external_connection.export
	);

	soc_system_command_e0 settings_acceleration_e0 (
		.clk        (clk_clk),                                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                          //               reset.reset_n
		.address    (mm_interconnect_1_settings_acceleration_e0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_settings_acceleration_e0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_settings_acceleration_e0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_settings_acceleration_e0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_settings_acceleration_e0_s1_readdata),   //                    .readdata
		.out_port   (settings_acceleration_e0_external_connection_export)       // external_connection.export
	);

	soc_system_command_e0 settings_acceleration_e1 (
		.clk        (clk_clk),                                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                          //               reset.reset_n
		.address    (mm_interconnect_1_settings_acceleration_e1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_settings_acceleration_e1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_settings_acceleration_e1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_settings_acceleration_e1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_settings_acceleration_e1_s1_readdata),   //                    .readdata
		.out_port   (settings_acceleration_e1_external_connection_export)       // external_connection.export
	);

	soc_system_command_e0 settings_acceleration_x (
		.clk        (clk_clk),                                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                         //               reset.reset_n
		.address    (mm_interconnect_1_settings_acceleration_x_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_settings_acceleration_x_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_settings_acceleration_x_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_settings_acceleration_x_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_settings_acceleration_x_s1_readdata),   //                    .readdata
		.out_port   (settings_acceleration_x_external_connection_export)       // external_connection.export
	);

	soc_system_command_e0 settings_acceleration_y (
		.clk        (clk_clk),                                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                         //               reset.reset_n
		.address    (mm_interconnect_1_settings_acceleration_y_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_settings_acceleration_y_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_settings_acceleration_y_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_settings_acceleration_y_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_settings_acceleration_y_s1_readdata),   //                    .readdata
		.out_port   (settings_acceleration_y_external_connection_export)       // external_connection.export
	);

	soc_system_command_e0 settings_acceleration_z (
		.clk        (clk_clk),                                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                         //               reset.reset_n
		.address    (mm_interconnect_1_settings_acceleration_z_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_settings_acceleration_z_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_settings_acceleration_z_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_settings_acceleration_z_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_settings_acceleration_z_s1_readdata),   //                    .readdata
		.out_port   (settings_acceleration_z_external_connection_export)       // external_connection.export
	);

	soc_system_command_e0 settings_jerk_e0 (
		.clk        (clk_clk),                                          //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                  //               reset.reset_n
		.address    (mm_interconnect_1_settings_jerk_e0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_settings_jerk_e0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_settings_jerk_e0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_settings_jerk_e0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_settings_jerk_e0_s1_readdata),   //                    .readdata
		.out_port   (settings_jerk_e0_external_connection_export)       // external_connection.export
	);

	soc_system_command_e0 settings_jerk_e1 (
		.clk        (clk_clk),                                          //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                  //               reset.reset_n
		.address    (mm_interconnect_1_settings_jerk_e1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_settings_jerk_e1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_settings_jerk_e1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_settings_jerk_e1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_settings_jerk_e1_s1_readdata),   //                    .readdata
		.out_port   (settings_jerk_e1_external_connection_export)       // external_connection.export
	);

	soc_system_command_e0 settings_jerk_x (
		.clk        (clk_clk),                                         //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                 //               reset.reset_n
		.address    (mm_interconnect_1_settings_jerk_x_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_settings_jerk_x_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_settings_jerk_x_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_settings_jerk_x_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_settings_jerk_x_s1_readdata),   //                    .readdata
		.out_port   (settings_jerk_x_external_connection_export)       // external_connection.export
	);

	soc_system_command_e0 settings_jerk_y (
		.clk        (clk_clk),                                         //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                 //               reset.reset_n
		.address    (mm_interconnect_1_settings_jerk_y_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_settings_jerk_y_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_settings_jerk_y_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_settings_jerk_y_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_settings_jerk_y_s1_readdata),   //                    .readdata
		.out_port   (settings_jerk_y_external_connection_export)       // external_connection.export
	);

	soc_system_command_e0 settings_jerk_z (
		.clk        (clk_clk),                                         //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                 //               reset.reset_n
		.address    (mm_interconnect_1_settings_jerk_z_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_settings_jerk_z_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_settings_jerk_z_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_settings_jerk_z_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_settings_jerk_z_s1_readdata),   //                    .readdata
		.out_port   (settings_jerk_z_external_connection_export)       // external_connection.export
	);

	soc_system_command_e0 settings_max_speed_e0 (
		.clk        (clk_clk),                                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                       //               reset.reset_n
		.address    (mm_interconnect_1_settings_max_speed_e0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_settings_max_speed_e0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_settings_max_speed_e0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_settings_max_speed_e0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_settings_max_speed_e0_s1_readdata),   //                    .readdata
		.out_port   (settings_max_speed_e0_external_connection_export)       // external_connection.export
	);

	soc_system_command_e0 settings_max_speed_e1 (
		.clk        (clk_clk),                                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                       //               reset.reset_n
		.address    (mm_interconnect_1_settings_max_speed_e1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_settings_max_speed_e1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_settings_max_speed_e1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_settings_max_speed_e1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_settings_max_speed_e1_s1_readdata),   //                    .readdata
		.out_port   (settings_max_speed_e1_external_connection_export)       // external_connection.export
	);

	soc_system_command_e0 settings_max_speed_x (
		.clk        (clk_clk),                                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                      //               reset.reset_n
		.address    (mm_interconnect_1_settings_max_speed_x_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_settings_max_speed_x_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_settings_max_speed_x_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_settings_max_speed_x_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_settings_max_speed_x_s1_readdata),   //                    .readdata
		.out_port   (settings_max_speed_x_external_connection_export)       // external_connection.export
	);

	soc_system_command_e0 settings_max_speed_y (
		.clk        (clk_clk),                                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                      //               reset.reset_n
		.address    (mm_interconnect_1_settings_max_speed_y_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_settings_max_speed_y_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_settings_max_speed_y_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_settings_max_speed_y_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_settings_max_speed_y_s1_readdata),   //                    .readdata
		.out_port   (settings_max_speed_y_external_connection_export)       // external_connection.export
	);

	soc_system_command_e0 settings_max_speed_z (
		.clk        (clk_clk),                                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                      //               reset.reset_n
		.address    (mm_interconnect_1_settings_max_speed_z_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_settings_max_speed_z_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_settings_max_speed_z_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_settings_max_speed_z_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_settings_max_speed_z_s1_readdata),   //                    .readdata
		.out_port   (settings_max_speed_z_external_connection_export)       // external_connection.export
	);

	soc_system_command_dt settings_max_temp_bed (
		.clk        (clk_clk),                                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                       //               reset.reset_n
		.address    (mm_interconnect_1_settings_max_temp_bed_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_settings_max_temp_bed_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_settings_max_temp_bed_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_settings_max_temp_bed_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_settings_max_temp_bed_s1_readdata),   //                    .readdata
		.out_port   (settings_max_temp_bed_external_connection_export)       // external_connection.export
	);

	soc_system_command_dt settings_max_temp_e0 (
		.clk        (clk_clk),                                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                      //               reset.reset_n
		.address    (mm_interconnect_1_settings_max_temp_e0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_settings_max_temp_e0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_settings_max_temp_e0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_settings_max_temp_e0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_settings_max_temp_e0_s1_readdata),   //                    .readdata
		.out_port   (settings_max_temp_e0_external_connection_export)       // external_connection.export
	);

	soc_system_command_dt settings_max_temp_e1 (
		.clk        (clk_clk),                                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                      //               reset.reset_n
		.address    (mm_interconnect_1_settings_max_temp_e1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_settings_max_temp_e1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_settings_max_temp_e1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_settings_max_temp_e1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_settings_max_temp_e1_s1_readdata),   //                    .readdata
		.out_port   (settings_max_temp_e1_external_connection_export)       // external_connection.export
	);

	soc_system_flags_in step_e0_now (
		.clk      (clk_clk),                                   //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address  (mm_interconnect_1_step_e0_now_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_step_e0_now_s1_readdata), //                    .readdata
		.in_port  (step_e0_now_external_connection_export)     // external_connection.export
	);

	soc_system_flags_in step_e1_now (
		.clk      (clk_clk),                                   //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address  (mm_interconnect_1_step_e1_now_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_step_e1_now_s1_readdata), //                    .readdata
		.in_port  (step_e1_now_external_connection_export)     // external_connection.export
	);

	soc_system_flags_in step_x_now (
		.clk      (clk_clk),                                  //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_1_step_x_now_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_step_x_now_s1_readdata), //                    .readdata
		.in_port  (step_x_now_external_connection_export)     // external_connection.export
	);

	soc_system_flags_in step_y_now (
		.clk      (clk_clk),                                  //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_1_step_y_now_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_step_y_now_s1_readdata), //                    .readdata
		.in_port  (step_y_now_external_connection_export)     // external_connection.export
	);

	soc_system_flags_in step_z_now (
		.clk      (clk_clk),                                  //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_1_step_z_now_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_step_z_now_s1_readdata), //                    .readdata
		.in_port  (step_z_now_external_connection_export)     // external_connection.export
	);

	soc_system_sysid_qsys sysid_qsys (
		.clock    (clk_clk),                                             //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                     //         reset.reset_n
		.readdata (mm_interconnect_1_sysid_qsys_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_1_sysid_qsys_control_slave_address)   //              .address
	);

	soc_system_position_e0 temp_0 (
		.clk      (clk_clk),                              //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address  (mm_interconnect_1_temp_0_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_temp_0_s1_readdata), //                    .readdata
		.in_port  (temp_0_external_connection_export)     // external_connection.export
	);

	soc_system_position_e0 temp_1 (
		.clk      (clk_clk),                              //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address  (mm_interconnect_1_temp_1_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_temp_1_s1_readdata), //                    .readdata
		.in_port  (temp_1_external_connection_export)     // external_connection.export
	);

	soc_system_position_e0 temp_2 (
		.clk      (clk_clk),                              //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address  (mm_interconnect_1_temp_2_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_temp_2_s1_readdata), //                    .readdata
		.in_port  (temp_2_external_connection_export)     // external_connection.export
	);

	soc_system_flags_in timing_e0_0 (
		.clk      (clk_clk),                                   //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address  (mm_interconnect_1_timing_e0_0_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_timing_e0_0_s1_readdata), //                    .readdata
		.in_port  (timing_e0_0_external_connection_export)     // external_connection.export
	);

	soc_system_flags_in timing_e0_1 (
		.clk      (clk_clk),                                   //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address  (mm_interconnect_1_timing_e0_1_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_timing_e0_1_s1_readdata), //                    .readdata
		.in_port  (timing_e0_1_external_connection_export)     // external_connection.export
	);

	soc_system_flags_in timing_e0_2 (
		.clk      (clk_clk),                                   //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address  (mm_interconnect_1_timing_e0_2_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_timing_e0_2_s1_readdata), //                    .readdata
		.in_port  (timing_e0_2_external_connection_export)     // external_connection.export
	);

	soc_system_flags_in timing_e0_3 (
		.clk      (clk_clk),                                   //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address  (mm_interconnect_1_timing_e0_3_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_timing_e0_3_s1_readdata), //                    .readdata
		.in_port  (timing_e0_3_external_connection_export)     // external_connection.export
	);

	soc_system_flags_in timing_e1_0 (
		.clk      (clk_clk),                                   //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address  (mm_interconnect_1_timing_e1_0_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_timing_e1_0_s1_readdata), //                    .readdata
		.in_port  (timing_e1_0_external_connection_export)     // external_connection.export
	);

	soc_system_flags_in timing_e1_1 (
		.clk      (clk_clk),                                   //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address  (mm_interconnect_1_timing_e1_1_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_timing_e1_1_s1_readdata), //                    .readdata
		.in_port  (timing_e1_1_external_connection_export)     // external_connection.export
	);

	soc_system_flags_in timing_e1_2 (
		.clk      (clk_clk),                                   //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address  (mm_interconnect_1_timing_e1_2_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_timing_e1_2_s1_readdata), //                    .readdata
		.in_port  (timing_e1_2_external_connection_export)     // external_connection.export
	);

	soc_system_flags_in timing_e1_3 (
		.clk      (clk_clk),                                   //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address  (mm_interconnect_1_timing_e1_3_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_timing_e1_3_s1_readdata), //                    .readdata
		.in_port  (timing_e1_3_external_connection_export)     // external_connection.export
	);

	soc_system_flags_in timing_x_0 (
		.clk      (clk_clk),                                  //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_1_timing_x_0_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_timing_x_0_s1_readdata), //                    .readdata
		.in_port  (timing_x_0_external_connection_export)     // external_connection.export
	);

	soc_system_flags_in timing_x_1 (
		.clk      (clk_clk),                                  //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_1_timing_x_1_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_timing_x_1_s1_readdata), //                    .readdata
		.in_port  (timing_x_1_external_connection_export)     // external_connection.export
	);

	soc_system_flags_in timing_x_2 (
		.clk      (clk_clk),                                  //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_1_timing_x_2_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_timing_x_2_s1_readdata), //                    .readdata
		.in_port  (timing_x_2_external_connection_export)     // external_connection.export
	);

	soc_system_flags_in timing_x_3 (
		.clk      (clk_clk),                                  //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_1_timing_x_3_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_timing_x_3_s1_readdata), //                    .readdata
		.in_port  (timing_x_3_external_connection_export)     // external_connection.export
	);

	soc_system_flags_in timing_y_0 (
		.clk      (clk_clk),                                  //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_1_timing_y_0_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_timing_y_0_s1_readdata), //                    .readdata
		.in_port  (timing_y_0_external_connection_export)     // external_connection.export
	);

	soc_system_flags_in timing_y_1 (
		.clk      (clk_clk),                                  //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_1_timing_y_1_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_timing_y_1_s1_readdata), //                    .readdata
		.in_port  (timing_y_1_external_connection_export)     // external_connection.export
	);

	soc_system_flags_in timing_y_2 (
		.clk      (clk_clk),                                  //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_1_timing_y_2_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_timing_y_2_s1_readdata), //                    .readdata
		.in_port  (timing_y_2_external_connection_export)     // external_connection.export
	);

	soc_system_flags_in timing_y_3 (
		.clk      (clk_clk),                                  //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_1_timing_y_3_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_timing_y_3_s1_readdata), //                    .readdata
		.in_port  (timing_y_3_external_connection_export)     // external_connection.export
	);

	soc_system_flags_in timing_z_0 (
		.clk      (clk_clk),                                  //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_1_timing_z_0_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_timing_z_0_s1_readdata), //                    .readdata
		.in_port  (timing_z_0_external_connection_export)     // external_connection.export
	);

	soc_system_flags_in timing_z_1 (
		.clk      (clk_clk),                                  //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_1_timing_z_1_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_timing_z_1_s1_readdata), //                    .readdata
		.in_port  (timing_z_1_external_connection_export)     // external_connection.export
	);

	soc_system_flags_in timing_z_2 (
		.clk      (clk_clk),                                  //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_1_timing_z_2_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_timing_z_2_s1_readdata), //                    .readdata
		.in_port  (timing_z_2_external_connection_export)     // external_connection.export
	);

	soc_system_flags_in timing_z_3 (
		.clk      (clk_clk),                                  //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_1_timing_z_3_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_timing_z_3_s1_readdata), //                    .readdata
		.in_port  (timing_z_3_external_connection_export)     // external_connection.export
	);

	soc_system_mm_interconnect_0 mm_interconnect_0 (
		.hps_0_h2f_lw_axi_master_awid                                        (hps_0_h2f_lw_axi_master_awid),                   //                                       hps_0_h2f_lw_axi_master.awid
		.hps_0_h2f_lw_axi_master_awaddr                                      (hps_0_h2f_lw_axi_master_awaddr),                 //                                                              .awaddr
		.hps_0_h2f_lw_axi_master_awlen                                       (hps_0_h2f_lw_axi_master_awlen),                  //                                                              .awlen
		.hps_0_h2f_lw_axi_master_awsize                                      (hps_0_h2f_lw_axi_master_awsize),                 //                                                              .awsize
		.hps_0_h2f_lw_axi_master_awburst                                     (hps_0_h2f_lw_axi_master_awburst),                //                                                              .awburst
		.hps_0_h2f_lw_axi_master_awlock                                      (hps_0_h2f_lw_axi_master_awlock),                 //                                                              .awlock
		.hps_0_h2f_lw_axi_master_awcache                                     (hps_0_h2f_lw_axi_master_awcache),                //                                                              .awcache
		.hps_0_h2f_lw_axi_master_awprot                                      (hps_0_h2f_lw_axi_master_awprot),                 //                                                              .awprot
		.hps_0_h2f_lw_axi_master_awvalid                                     (hps_0_h2f_lw_axi_master_awvalid),                //                                                              .awvalid
		.hps_0_h2f_lw_axi_master_awready                                     (hps_0_h2f_lw_axi_master_awready),                //                                                              .awready
		.hps_0_h2f_lw_axi_master_wid                                         (hps_0_h2f_lw_axi_master_wid),                    //                                                              .wid
		.hps_0_h2f_lw_axi_master_wdata                                       (hps_0_h2f_lw_axi_master_wdata),                  //                                                              .wdata
		.hps_0_h2f_lw_axi_master_wstrb                                       (hps_0_h2f_lw_axi_master_wstrb),                  //                                                              .wstrb
		.hps_0_h2f_lw_axi_master_wlast                                       (hps_0_h2f_lw_axi_master_wlast),                  //                                                              .wlast
		.hps_0_h2f_lw_axi_master_wvalid                                      (hps_0_h2f_lw_axi_master_wvalid),                 //                                                              .wvalid
		.hps_0_h2f_lw_axi_master_wready                                      (hps_0_h2f_lw_axi_master_wready),                 //                                                              .wready
		.hps_0_h2f_lw_axi_master_bid                                         (hps_0_h2f_lw_axi_master_bid),                    //                                                              .bid
		.hps_0_h2f_lw_axi_master_bresp                                       (hps_0_h2f_lw_axi_master_bresp),                  //                                                              .bresp
		.hps_0_h2f_lw_axi_master_bvalid                                      (hps_0_h2f_lw_axi_master_bvalid),                 //                                                              .bvalid
		.hps_0_h2f_lw_axi_master_bready                                      (hps_0_h2f_lw_axi_master_bready),                 //                                                              .bready
		.hps_0_h2f_lw_axi_master_arid                                        (hps_0_h2f_lw_axi_master_arid),                   //                                                              .arid
		.hps_0_h2f_lw_axi_master_araddr                                      (hps_0_h2f_lw_axi_master_araddr),                 //                                                              .araddr
		.hps_0_h2f_lw_axi_master_arlen                                       (hps_0_h2f_lw_axi_master_arlen),                  //                                                              .arlen
		.hps_0_h2f_lw_axi_master_arsize                                      (hps_0_h2f_lw_axi_master_arsize),                 //                                                              .arsize
		.hps_0_h2f_lw_axi_master_arburst                                     (hps_0_h2f_lw_axi_master_arburst),                //                                                              .arburst
		.hps_0_h2f_lw_axi_master_arlock                                      (hps_0_h2f_lw_axi_master_arlock),                 //                                                              .arlock
		.hps_0_h2f_lw_axi_master_arcache                                     (hps_0_h2f_lw_axi_master_arcache),                //                                                              .arcache
		.hps_0_h2f_lw_axi_master_arprot                                      (hps_0_h2f_lw_axi_master_arprot),                 //                                                              .arprot
		.hps_0_h2f_lw_axi_master_arvalid                                     (hps_0_h2f_lw_axi_master_arvalid),                //                                                              .arvalid
		.hps_0_h2f_lw_axi_master_arready                                     (hps_0_h2f_lw_axi_master_arready),                //                                                              .arready
		.hps_0_h2f_lw_axi_master_rid                                         (hps_0_h2f_lw_axi_master_rid),                    //                                                              .rid
		.hps_0_h2f_lw_axi_master_rdata                                       (hps_0_h2f_lw_axi_master_rdata),                  //                                                              .rdata
		.hps_0_h2f_lw_axi_master_rresp                                       (hps_0_h2f_lw_axi_master_rresp),                  //                                                              .rresp
		.hps_0_h2f_lw_axi_master_rlast                                       (hps_0_h2f_lw_axi_master_rlast),                  //                                                              .rlast
		.hps_0_h2f_lw_axi_master_rvalid                                      (hps_0_h2f_lw_axi_master_rvalid),                 //                                                              .rvalid
		.hps_0_h2f_lw_axi_master_rready                                      (hps_0_h2f_lw_axi_master_rready),                 //                                                              .rready
		.clk_0_clk_clk                                                       (clk_clk),                                        //                                                     clk_0_clk.clk
		.hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),             // hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.mm_bridge_0_reset_reset_bridge_in_reset_reset                       (rst_controller_reset_out_reset),                 //                       mm_bridge_0_reset_reset_bridge_in_reset.reset
		.mm_bridge_0_s0_address                                              (mm_interconnect_0_mm_bridge_0_s0_address),       //                                                mm_bridge_0_s0.address
		.mm_bridge_0_s0_write                                                (mm_interconnect_0_mm_bridge_0_s0_write),         //                                                              .write
		.mm_bridge_0_s0_read                                                 (mm_interconnect_0_mm_bridge_0_s0_read),          //                                                              .read
		.mm_bridge_0_s0_readdata                                             (mm_interconnect_0_mm_bridge_0_s0_readdata),      //                                                              .readdata
		.mm_bridge_0_s0_writedata                                            (mm_interconnect_0_mm_bridge_0_s0_writedata),     //                                                              .writedata
		.mm_bridge_0_s0_burstcount                                           (mm_interconnect_0_mm_bridge_0_s0_burstcount),    //                                                              .burstcount
		.mm_bridge_0_s0_byteenable                                           (mm_interconnect_0_mm_bridge_0_s0_byteenable),    //                                                              .byteenable
		.mm_bridge_0_s0_readdatavalid                                        (mm_interconnect_0_mm_bridge_0_s0_readdatavalid), //                                                              .readdatavalid
		.mm_bridge_0_s0_waitrequest                                          (mm_interconnect_0_mm_bridge_0_s0_waitrequest),   //                                                              .waitrequest
		.mm_bridge_0_s0_debugaccess                                          (mm_interconnect_0_mm_bridge_0_s0_debugaccess)    //                                                              .debugaccess
	);

	soc_system_mm_interconnect_1 mm_interconnect_1 (
		.clk_0_clk_clk                                          (clk_clk),                                                   //                                        clk_0_clk.clk
		.fpga_only_master_clk_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                            // fpga_only_master_clk_reset_reset_bridge_in_reset.reset
		.mm_bridge_0_reset_reset_bridge_in_reset_reset          (rst_controller_reset_out_reset),                            //          mm_bridge_0_reset_reset_bridge_in_reset.reset
		.fpga_only_master_master_address                        (fpga_only_master_master_address),                           //                          fpga_only_master_master.address
		.fpga_only_master_master_waitrequest                    (fpga_only_master_master_waitrequest),                       //                                                 .waitrequest
		.fpga_only_master_master_byteenable                     (fpga_only_master_master_byteenable),                        //                                                 .byteenable
		.fpga_only_master_master_read                           (fpga_only_master_master_read),                              //                                                 .read
		.fpga_only_master_master_readdata                       (fpga_only_master_master_readdata),                          //                                                 .readdata
		.fpga_only_master_master_readdatavalid                  (fpga_only_master_master_readdatavalid),                     //                                                 .readdatavalid
		.fpga_only_master_master_write                          (fpga_only_master_master_write),                             //                                                 .write
		.fpga_only_master_master_writedata                      (fpga_only_master_master_writedata),                         //                                                 .writedata
		.mm_bridge_0_m0_address                                 (mm_bridge_0_m0_address),                                    //                                   mm_bridge_0_m0.address
		.mm_bridge_0_m0_waitrequest                             (mm_bridge_0_m0_waitrequest),                                //                                                 .waitrequest
		.mm_bridge_0_m0_burstcount                              (mm_bridge_0_m0_burstcount),                                 //                                                 .burstcount
		.mm_bridge_0_m0_byteenable                              (mm_bridge_0_m0_byteenable),                                 //                                                 .byteenable
		.mm_bridge_0_m0_read                                    (mm_bridge_0_m0_read),                                       //                                                 .read
		.mm_bridge_0_m0_readdata                                (mm_bridge_0_m0_readdata),                                   //                                                 .readdata
		.mm_bridge_0_m0_readdatavalid                           (mm_bridge_0_m0_readdatavalid),                              //                                                 .readdatavalid
		.mm_bridge_0_m0_write                                   (mm_bridge_0_m0_write),                                      //                                                 .write
		.mm_bridge_0_m0_writedata                               (mm_bridge_0_m0_writedata),                                  //                                                 .writedata
		.mm_bridge_0_m0_debugaccess                             (mm_bridge_0_m0_debugaccess),                                //                                                 .debugaccess
		.command_dt_s1_address                                  (mm_interconnect_1_command_dt_s1_address),                   //                                    command_dt_s1.address
		.command_dt_s1_write                                    (mm_interconnect_1_command_dt_s1_write),                     //                                                 .write
		.command_dt_s1_readdata                                 (mm_interconnect_1_command_dt_s1_readdata),                  //                                                 .readdata
		.command_dt_s1_writedata                                (mm_interconnect_1_command_dt_s1_writedata),                 //                                                 .writedata
		.command_dt_s1_chipselect                               (mm_interconnect_1_command_dt_s1_chipselect),                //                                                 .chipselect
		.command_e0_s1_address                                  (mm_interconnect_1_command_e0_s1_address),                   //                                    command_e0_s1.address
		.command_e0_s1_write                                    (mm_interconnect_1_command_e0_s1_write),                     //                                                 .write
		.command_e0_s1_readdata                                 (mm_interconnect_1_command_e0_s1_readdata),                  //                                                 .readdata
		.command_e0_s1_writedata                                (mm_interconnect_1_command_e0_s1_writedata),                 //                                                 .writedata
		.command_e0_s1_chipselect                               (mm_interconnect_1_command_e0_s1_chipselect),                //                                                 .chipselect
		.command_e1_s1_address                                  (mm_interconnect_1_command_e1_s1_address),                   //                                    command_e1_s1.address
		.command_e1_s1_write                                    (mm_interconnect_1_command_e1_s1_write),                     //                                                 .write
		.command_e1_s1_readdata                                 (mm_interconnect_1_command_e1_s1_readdata),                  //                                                 .readdata
		.command_e1_s1_writedata                                (mm_interconnect_1_command_e1_s1_writedata),                 //                                                 .writedata
		.command_e1_s1_chipselect                               (mm_interconnect_1_command_e1_s1_chipselect),                //                                                 .chipselect
		.command_f_e0_s1_address                                (mm_interconnect_1_command_f_e0_s1_address),                 //                                  command_f_e0_s1.address
		.command_f_e0_s1_write                                  (mm_interconnect_1_command_f_e0_s1_write),                   //                                                 .write
		.command_f_e0_s1_readdata                               (mm_interconnect_1_command_f_e0_s1_readdata),                //                                                 .readdata
		.command_f_e0_s1_writedata                              (mm_interconnect_1_command_f_e0_s1_writedata),               //                                                 .writedata
		.command_f_e0_s1_chipselect                             (mm_interconnect_1_command_f_e0_s1_chipselect),              //                                                 .chipselect
		.command_f_e1_s1_address                                (mm_interconnect_1_command_f_e1_s1_address),                 //                                  command_f_e1_s1.address
		.command_f_e1_s1_write                                  (mm_interconnect_1_command_f_e1_s1_write),                   //                                                 .write
		.command_f_e1_s1_readdata                               (mm_interconnect_1_command_f_e1_s1_readdata),                //                                                 .readdata
		.command_f_e1_s1_writedata                              (mm_interconnect_1_command_f_e1_s1_writedata),               //                                                 .writedata
		.command_f_e1_s1_chipselect                             (mm_interconnect_1_command_f_e1_s1_chipselect),              //                                                 .chipselect
		.command_f_x_s1_address                                 (mm_interconnect_1_command_f_x_s1_address),                  //                                   command_f_x_s1.address
		.command_f_x_s1_write                                   (mm_interconnect_1_command_f_x_s1_write),                    //                                                 .write
		.command_f_x_s1_readdata                                (mm_interconnect_1_command_f_x_s1_readdata),                 //                                                 .readdata
		.command_f_x_s1_writedata                               (mm_interconnect_1_command_f_x_s1_writedata),                //                                                 .writedata
		.command_f_x_s1_chipselect                              (mm_interconnect_1_command_f_x_s1_chipselect),               //                                                 .chipselect
		.command_f_y_s1_address                                 (mm_interconnect_1_command_f_y_s1_address),                  //                                   command_f_y_s1.address
		.command_f_y_s1_write                                   (mm_interconnect_1_command_f_y_s1_write),                    //                                                 .write
		.command_f_y_s1_readdata                                (mm_interconnect_1_command_f_y_s1_readdata),                 //                                                 .readdata
		.command_f_y_s1_writedata                               (mm_interconnect_1_command_f_y_s1_writedata),                //                                                 .writedata
		.command_f_y_s1_chipselect                              (mm_interconnect_1_command_f_y_s1_chipselect),               //                                                 .chipselect
		.command_f_z_s1_address                                 (mm_interconnect_1_command_f_z_s1_address),                  //                                   command_f_z_s1.address
		.command_f_z_s1_write                                   (mm_interconnect_1_command_f_z_s1_write),                    //                                                 .write
		.command_f_z_s1_readdata                                (mm_interconnect_1_command_f_z_s1_readdata),                 //                                                 .readdata
		.command_f_z_s1_writedata                               (mm_interconnect_1_command_f_z_s1_writedata),                //                                                 .writedata
		.command_f_z_s1_chipselect                              (mm_interconnect_1_command_f_z_s1_chipselect),               //                                                 .chipselect
		.command_t_s1_address                                   (mm_interconnect_1_command_t_s1_address),                    //                                     command_t_s1.address
		.command_t_s1_write                                     (mm_interconnect_1_command_t_s1_write),                      //                                                 .write
		.command_t_s1_readdata                                  (mm_interconnect_1_command_t_s1_readdata),                   //                                                 .readdata
		.command_t_s1_writedata                                 (mm_interconnect_1_command_t_s1_writedata),                  //                                                 .writedata
		.command_t_s1_chipselect                                (mm_interconnect_1_command_t_s1_chipselect),                 //                                                 .chipselect
		.command_type_s1_address                                (mm_interconnect_1_command_type_s1_address),                 //                                  command_type_s1.address
		.command_type_s1_write                                  (mm_interconnect_1_command_type_s1_write),                   //                                                 .write
		.command_type_s1_readdata                               (mm_interconnect_1_command_type_s1_readdata),                //                                                 .readdata
		.command_type_s1_writedata                              (mm_interconnect_1_command_type_s1_writedata),               //                                                 .writedata
		.command_type_s1_chipselect                             (mm_interconnect_1_command_type_s1_chipselect),              //                                                 .chipselect
		.command_x_s1_address                                   (mm_interconnect_1_command_x_s1_address),                    //                                     command_x_s1.address
		.command_x_s1_write                                     (mm_interconnect_1_command_x_s1_write),                      //                                                 .write
		.command_x_s1_readdata                                  (mm_interconnect_1_command_x_s1_readdata),                   //                                                 .readdata
		.command_x_s1_writedata                                 (mm_interconnect_1_command_x_s1_writedata),                  //                                                 .writedata
		.command_x_s1_chipselect                                (mm_interconnect_1_command_x_s1_chipselect),                 //                                                 .chipselect
		.command_y_s1_address                                   (mm_interconnect_1_command_y_s1_address),                    //                                     command_y_s1.address
		.command_y_s1_write                                     (mm_interconnect_1_command_y_s1_write),                      //                                                 .write
		.command_y_s1_readdata                                  (mm_interconnect_1_command_y_s1_readdata),                   //                                                 .readdata
		.command_y_s1_writedata                                 (mm_interconnect_1_command_y_s1_writedata),                  //                                                 .writedata
		.command_y_s1_chipselect                                (mm_interconnect_1_command_y_s1_chipselect),                 //                                                 .chipselect
		.command_z_s1_address                                   (mm_interconnect_1_command_z_s1_address),                    //                                     command_z_s1.address
		.command_z_s1_write                                     (mm_interconnect_1_command_z_s1_write),                      //                                                 .write
		.command_z_s1_readdata                                  (mm_interconnect_1_command_z_s1_readdata),                   //                                                 .readdata
		.command_z_s1_writedata                                 (mm_interconnect_1_command_z_s1_writedata),                  //                                                 .writedata
		.command_z_s1_chipselect                                (mm_interconnect_1_command_z_s1_chipselect),                 //                                                 .chipselect
		.flags_in_s1_address                                    (mm_interconnect_1_flags_in_s1_address),                     //                                      flags_in_s1.address
		.flags_in_s1_readdata                                   (mm_interconnect_1_flags_in_s1_readdata),                    //                                                 .readdata
		.flags_out_s1_address                                   (mm_interconnect_1_flags_out_s1_address),                    //                                     flags_out_s1.address
		.flags_out_s1_write                                     (mm_interconnect_1_flags_out_s1_write),                      //                                                 .write
		.flags_out_s1_readdata                                  (mm_interconnect_1_flags_out_s1_readdata),                   //                                                 .readdata
		.flags_out_s1_writedata                                 (mm_interconnect_1_flags_out_s1_writedata),                  //                                                 .writedata
		.flags_out_s1_chipselect                                (mm_interconnect_1_flags_out_s1_chipselect),                 //                                                 .chipselect
		.ILC_avalon_slave_address                               (mm_interconnect_1_ilc_avalon_slave_address),                //                                 ILC_avalon_slave.address
		.ILC_avalon_slave_write                                 (mm_interconnect_1_ilc_avalon_slave_write),                  //                                                 .write
		.ILC_avalon_slave_read                                  (mm_interconnect_1_ilc_avalon_slave_read),                   //                                                 .read
		.ILC_avalon_slave_readdata                              (mm_interconnect_1_ilc_avalon_slave_readdata),               //                                                 .readdata
		.ILC_avalon_slave_writedata                             (mm_interconnect_1_ilc_avalon_slave_writedata),              //                                                 .writedata
		.jtag_uart_avalon_jtag_slave_address                    (mm_interconnect_1_jtag_uart_avalon_jtag_slave_address),     //                      jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                      (mm_interconnect_1_jtag_uart_avalon_jtag_slave_write),       //                                                 .write
		.jtag_uart_avalon_jtag_slave_read                       (mm_interconnect_1_jtag_uart_avalon_jtag_slave_read),        //                                                 .read
		.jtag_uart_avalon_jtag_slave_readdata                   (mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata),    //                                                 .readdata
		.jtag_uart_avalon_jtag_slave_writedata                  (mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata),   //                                                 .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest                (mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest), //                                                 .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect                 (mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect),  //                                                 .chipselect
		.max_params_0_s1_address                                (mm_interconnect_1_max_params_0_s1_address),                 //                                  max_params_0_s1.address
		.max_params_0_s1_readdata                               (mm_interconnect_1_max_params_0_s1_readdata),                //                                                 .readdata
		.max_params_1_s1_address                                (mm_interconnect_1_max_params_1_s1_address),                 //                                  max_params_1_s1.address
		.max_params_1_s1_readdata                               (mm_interconnect_1_max_params_1_s1_readdata),                //                                                 .readdata
		.max_params_2_s1_address                                (mm_interconnect_1_max_params_2_s1_address),                 //                                  max_params_2_s1.address
		.max_params_2_s1_readdata                               (mm_interconnect_1_max_params_2_s1_readdata),                //                                                 .readdata
		.max_params_3_s1_address                                (mm_interconnect_1_max_params_3_s1_address),                 //                                  max_params_3_s1.address
		.max_params_3_s1_readdata                               (mm_interconnect_1_max_params_3_s1_readdata),                //                                                 .readdata
		.max_params_4_s1_address                                (mm_interconnect_1_max_params_4_s1_address),                 //                                  max_params_4_s1.address
		.max_params_4_s1_readdata                               (mm_interconnect_1_max_params_4_s1_readdata),                //                                                 .readdata
		.max_timing_0_s1_address                                (mm_interconnect_1_max_timing_0_s1_address),                 //                                  max_timing_0_s1.address
		.max_timing_0_s1_readdata                               (mm_interconnect_1_max_timing_0_s1_readdata),                //                                                 .readdata
		.max_timing_1_s1_address                                (mm_interconnect_1_max_timing_1_s1_address),                 //                                  max_timing_1_s1.address
		.max_timing_1_s1_readdata                               (mm_interconnect_1_max_timing_1_s1_readdata),                //                                                 .readdata
		.max_timing_2_s1_address                                (mm_interconnect_1_max_timing_2_s1_address),                 //                                  max_timing_2_s1.address
		.max_timing_2_s1_readdata                               (mm_interconnect_1_max_timing_2_s1_readdata),                //                                                 .readdata
		.max_timing_3_s1_address                                (mm_interconnect_1_max_timing_3_s1_address),                 //                                  max_timing_3_s1.address
		.max_timing_3_s1_readdata                               (mm_interconnect_1_max_timing_3_s1_readdata),                //                                                 .readdata
		.new_rparams_e0_0_s1_address                            (mm_interconnect_1_new_rparams_e0_0_s1_address),             //                              new_rparams_e0_0_s1.address
		.new_rparams_e0_0_s1_readdata                           (mm_interconnect_1_new_rparams_e0_0_s1_readdata),            //                                                 .readdata
		.new_rparams_e0_1_s1_address                            (mm_interconnect_1_new_rparams_e0_1_s1_address),             //                              new_rparams_e0_1_s1.address
		.new_rparams_e0_1_s1_readdata                           (mm_interconnect_1_new_rparams_e0_1_s1_readdata),            //                                                 .readdata
		.new_rparams_e0_2_s1_address                            (mm_interconnect_1_new_rparams_e0_2_s1_address),             //                              new_rparams_e0_2_s1.address
		.new_rparams_e0_2_s1_readdata                           (mm_interconnect_1_new_rparams_e0_2_s1_readdata),            //                                                 .readdata
		.new_rparams_e0_3_s1_address                            (mm_interconnect_1_new_rparams_e0_3_s1_address),             //                              new_rparams_e0_3_s1.address
		.new_rparams_e0_3_s1_readdata                           (mm_interconnect_1_new_rparams_e0_3_s1_readdata),            //                                                 .readdata
		.new_rparams_e0_4_s1_address                            (mm_interconnect_1_new_rparams_e0_4_s1_address),             //                              new_rparams_e0_4_s1.address
		.new_rparams_e0_4_s1_readdata                           (mm_interconnect_1_new_rparams_e0_4_s1_readdata),            //                                                 .readdata
		.new_rparams_e1_0_s1_address                            (mm_interconnect_1_new_rparams_e1_0_s1_address),             //                              new_rparams_e1_0_s1.address
		.new_rparams_e1_0_s1_readdata                           (mm_interconnect_1_new_rparams_e1_0_s1_readdata),            //                                                 .readdata
		.new_rparams_e1_1_s1_address                            (mm_interconnect_1_new_rparams_e1_1_s1_address),             //                              new_rparams_e1_1_s1.address
		.new_rparams_e1_1_s1_readdata                           (mm_interconnect_1_new_rparams_e1_1_s1_readdata),            //                                                 .readdata
		.new_rparams_e1_2_s1_address                            (mm_interconnect_1_new_rparams_e1_2_s1_address),             //                              new_rparams_e1_2_s1.address
		.new_rparams_e1_2_s1_readdata                           (mm_interconnect_1_new_rparams_e1_2_s1_readdata),            //                                                 .readdata
		.new_rparams_e1_3_s1_address                            (mm_interconnect_1_new_rparams_e1_3_s1_address),             //                              new_rparams_e1_3_s1.address
		.new_rparams_e1_3_s1_readdata                           (mm_interconnect_1_new_rparams_e1_3_s1_readdata),            //                                                 .readdata
		.new_rparams_e1_4_s1_address                            (mm_interconnect_1_new_rparams_e1_4_s1_address),             //                              new_rparams_e1_4_s1.address
		.new_rparams_e1_4_s1_readdata                           (mm_interconnect_1_new_rparams_e1_4_s1_readdata),            //                                                 .readdata
		.new_rparams_x_0_s1_address                             (mm_interconnect_1_new_rparams_x_0_s1_address),              //                               new_rparams_x_0_s1.address
		.new_rparams_x_0_s1_readdata                            (mm_interconnect_1_new_rparams_x_0_s1_readdata),             //                                                 .readdata
		.new_rparams_x_1_s1_address                             (mm_interconnect_1_new_rparams_x_1_s1_address),              //                               new_rparams_x_1_s1.address
		.new_rparams_x_1_s1_readdata                            (mm_interconnect_1_new_rparams_x_1_s1_readdata),             //                                                 .readdata
		.new_rparams_x_2_s1_address                             (mm_interconnect_1_new_rparams_x_2_s1_address),              //                               new_rparams_x_2_s1.address
		.new_rparams_x_2_s1_readdata                            (mm_interconnect_1_new_rparams_x_2_s1_readdata),             //                                                 .readdata
		.new_rparams_x_3_s1_address                             (mm_interconnect_1_new_rparams_x_3_s1_address),              //                               new_rparams_x_3_s1.address
		.new_rparams_x_3_s1_readdata                            (mm_interconnect_1_new_rparams_x_3_s1_readdata),             //                                                 .readdata
		.new_rparams_x_4_s1_address                             (mm_interconnect_1_new_rparams_x_4_s1_address),              //                               new_rparams_x_4_s1.address
		.new_rparams_x_4_s1_readdata                            (mm_interconnect_1_new_rparams_x_4_s1_readdata),             //                                                 .readdata
		.new_rparams_y_0_s1_address                             (mm_interconnect_1_new_rparams_y_0_s1_address),              //                               new_rparams_y_0_s1.address
		.new_rparams_y_0_s1_readdata                            (mm_interconnect_1_new_rparams_y_0_s1_readdata),             //                                                 .readdata
		.new_rparams_y_1_s1_address                             (mm_interconnect_1_new_rparams_y_1_s1_address),              //                               new_rparams_y_1_s1.address
		.new_rparams_y_1_s1_readdata                            (mm_interconnect_1_new_rparams_y_1_s1_readdata),             //                                                 .readdata
		.new_rparams_y_2_s1_address                             (mm_interconnect_1_new_rparams_y_2_s1_address),              //                               new_rparams_y_2_s1.address
		.new_rparams_y_2_s1_readdata                            (mm_interconnect_1_new_rparams_y_2_s1_readdata),             //                                                 .readdata
		.new_rparams_y_3_s1_address                             (mm_interconnect_1_new_rparams_y_3_s1_address),              //                               new_rparams_y_3_s1.address
		.new_rparams_y_3_s1_readdata                            (mm_interconnect_1_new_rparams_y_3_s1_readdata),             //                                                 .readdata
		.new_rparams_y_4_s1_address                             (mm_interconnect_1_new_rparams_y_4_s1_address),              //                               new_rparams_y_4_s1.address
		.new_rparams_y_4_s1_readdata                            (mm_interconnect_1_new_rparams_y_4_s1_readdata),             //                                                 .readdata
		.new_rparams_z_0_s1_address                             (mm_interconnect_1_new_rparams_z_0_s1_address),              //                               new_rparams_z_0_s1.address
		.new_rparams_z_0_s1_readdata                            (mm_interconnect_1_new_rparams_z_0_s1_readdata),             //                                                 .readdata
		.new_rparams_z_1_s1_address                             (mm_interconnect_1_new_rparams_z_1_s1_address),              //                               new_rparams_z_1_s1.address
		.new_rparams_z_1_s1_readdata                            (mm_interconnect_1_new_rparams_z_1_s1_readdata),             //                                                 .readdata
		.new_rparams_z_2_s1_address                             (mm_interconnect_1_new_rparams_z_2_s1_address),              //                               new_rparams_z_2_s1.address
		.new_rparams_z_2_s1_readdata                            (mm_interconnect_1_new_rparams_z_2_s1_readdata),             //                                                 .readdata
		.new_rparams_z_3_s1_address                             (mm_interconnect_1_new_rparams_z_3_s1_address),              //                               new_rparams_z_3_s1.address
		.new_rparams_z_3_s1_readdata                            (mm_interconnect_1_new_rparams_z_3_s1_readdata),             //                                                 .readdata
		.new_rparams_z_4_s1_address                             (mm_interconnect_1_new_rparams_z_4_s1_address),              //                               new_rparams_z_4_s1.address
		.new_rparams_z_4_s1_readdata                            (mm_interconnect_1_new_rparams_z_4_s1_readdata),             //                                                 .readdata
		.params_e0_0_s1_address                                 (mm_interconnect_1_params_e0_0_s1_address),                  //                                   params_e0_0_s1.address
		.params_e0_0_s1_readdata                                (mm_interconnect_1_params_e0_0_s1_readdata),                 //                                                 .readdata
		.params_e0_1_s1_address                                 (mm_interconnect_1_params_e0_1_s1_address),                  //                                   params_e0_1_s1.address
		.params_e0_1_s1_readdata                                (mm_interconnect_1_params_e0_1_s1_readdata),                 //                                                 .readdata
		.params_e0_2_s1_address                                 (mm_interconnect_1_params_e0_2_s1_address),                  //                                   params_e0_2_s1.address
		.params_e0_2_s1_readdata                                (mm_interconnect_1_params_e0_2_s1_readdata),                 //                                                 .readdata
		.params_e0_3_s1_address                                 (mm_interconnect_1_params_e0_3_s1_address),                  //                                   params_e0_3_s1.address
		.params_e0_3_s1_readdata                                (mm_interconnect_1_params_e0_3_s1_readdata),                 //                                                 .readdata
		.params_e0_4_s1_address                                 (mm_interconnect_1_params_e0_4_s1_address),                  //                                   params_e0_4_s1.address
		.params_e0_4_s1_readdata                                (mm_interconnect_1_params_e0_4_s1_readdata),                 //                                                 .readdata
		.params_e1_0_s1_address                                 (mm_interconnect_1_params_e1_0_s1_address),                  //                                   params_e1_0_s1.address
		.params_e1_0_s1_readdata                                (mm_interconnect_1_params_e1_0_s1_readdata),                 //                                                 .readdata
		.params_e1_1_s1_address                                 (mm_interconnect_1_params_e1_1_s1_address),                  //                                   params_e1_1_s1.address
		.params_e1_1_s1_readdata                                (mm_interconnect_1_params_e1_1_s1_readdata),                 //                                                 .readdata
		.params_e1_2_s1_address                                 (mm_interconnect_1_params_e1_2_s1_address),                  //                                   params_e1_2_s1.address
		.params_e1_2_s1_readdata                                (mm_interconnect_1_params_e1_2_s1_readdata),                 //                                                 .readdata
		.params_e1_3_s1_address                                 (mm_interconnect_1_params_e1_3_s1_address),                  //                                   params_e1_3_s1.address
		.params_e1_3_s1_readdata                                (mm_interconnect_1_params_e1_3_s1_readdata),                 //                                                 .readdata
		.params_e1_4_s1_address                                 (mm_interconnect_1_params_e1_4_s1_address),                  //                                   params_e1_4_s1.address
		.params_e1_4_s1_readdata                                (mm_interconnect_1_params_e1_4_s1_readdata),                 //                                                 .readdata
		.params_x_0_s1_address                                  (mm_interconnect_1_params_x_0_s1_address),                   //                                    params_x_0_s1.address
		.params_x_0_s1_readdata                                 (mm_interconnect_1_params_x_0_s1_readdata),                  //                                                 .readdata
		.params_x_1_s1_address                                  (mm_interconnect_1_params_x_1_s1_address),                   //                                    params_x_1_s1.address
		.params_x_1_s1_readdata                                 (mm_interconnect_1_params_x_1_s1_readdata),                  //                                                 .readdata
		.params_x_2_s1_address                                  (mm_interconnect_1_params_x_2_s1_address),                   //                                    params_x_2_s1.address
		.params_x_2_s1_readdata                                 (mm_interconnect_1_params_x_2_s1_readdata),                  //                                                 .readdata
		.params_x_3_s1_address                                  (mm_interconnect_1_params_x_3_s1_address),                   //                                    params_x_3_s1.address
		.params_x_3_s1_readdata                                 (mm_interconnect_1_params_x_3_s1_readdata),                  //                                                 .readdata
		.params_x_4_s1_address                                  (mm_interconnect_1_params_x_4_s1_address),                   //                                    params_x_4_s1.address
		.params_x_4_s1_readdata                                 (mm_interconnect_1_params_x_4_s1_readdata),                  //                                                 .readdata
		.params_y_0_s1_address                                  (mm_interconnect_1_params_y_0_s1_address),                   //                                    params_y_0_s1.address
		.params_y_0_s1_readdata                                 (mm_interconnect_1_params_y_0_s1_readdata),                  //                                                 .readdata
		.params_y_1_s1_address                                  (mm_interconnect_1_params_y_1_s1_address),                   //                                    params_y_1_s1.address
		.params_y_1_s1_readdata                                 (mm_interconnect_1_params_y_1_s1_readdata),                  //                                                 .readdata
		.params_y_2_s1_address                                  (mm_interconnect_1_params_y_2_s1_address),                   //                                    params_y_2_s1.address
		.params_y_2_s1_readdata                                 (mm_interconnect_1_params_y_2_s1_readdata),                  //                                                 .readdata
		.params_y_3_s1_address                                  (mm_interconnect_1_params_y_3_s1_address),                   //                                    params_y_3_s1.address
		.params_y_3_s1_readdata                                 (mm_interconnect_1_params_y_3_s1_readdata),                  //                                                 .readdata
		.params_y_4_s1_address                                  (mm_interconnect_1_params_y_4_s1_address),                   //                                    params_y_4_s1.address
		.params_y_4_s1_readdata                                 (mm_interconnect_1_params_y_4_s1_readdata),                  //                                                 .readdata
		.params_z_0_s1_address                                  (mm_interconnect_1_params_z_0_s1_address),                   //                                    params_z_0_s1.address
		.params_z_0_s1_readdata                                 (mm_interconnect_1_params_z_0_s1_readdata),                  //                                                 .readdata
		.params_z_1_s1_address                                  (mm_interconnect_1_params_z_1_s1_address),                   //                                    params_z_1_s1.address
		.params_z_1_s1_readdata                                 (mm_interconnect_1_params_z_1_s1_readdata),                  //                                                 .readdata
		.params_z_2_s1_address                                  (mm_interconnect_1_params_z_2_s1_address),                   //                                    params_z_2_s1.address
		.params_z_2_s1_readdata                                 (mm_interconnect_1_params_z_2_s1_readdata),                  //                                                 .readdata
		.params_z_3_s1_address                                  (mm_interconnect_1_params_z_3_s1_address),                   //                                    params_z_3_s1.address
		.params_z_3_s1_readdata                                 (mm_interconnect_1_params_z_3_s1_readdata),                  //                                                 .readdata
		.params_z_4_s1_address                                  (mm_interconnect_1_params_z_4_s1_address),                   //                                    params_z_4_s1.address
		.params_z_4_s1_readdata                                 (mm_interconnect_1_params_z_4_s1_readdata),                  //                                                 .readdata
		.position_e0_s1_address                                 (mm_interconnect_1_position_e0_s1_address),                  //                                   position_e0_s1.address
		.position_e0_s1_readdata                                (mm_interconnect_1_position_e0_s1_readdata),                 //                                                 .readdata
		.position_e1_s1_address                                 (mm_interconnect_1_position_e1_s1_address),                  //                                   position_e1_s1.address
		.position_e1_s1_readdata                                (mm_interconnect_1_position_e1_s1_readdata),                 //                                                 .readdata
		.position_x_s1_address                                  (mm_interconnect_1_position_x_s1_address),                   //                                    position_x_s1.address
		.position_x_s1_readdata                                 (mm_interconnect_1_position_x_s1_readdata),                  //                                                 .readdata
		.position_y_s1_address                                  (mm_interconnect_1_position_y_s1_address),                   //                                    position_y_s1.address
		.position_y_s1_readdata                                 (mm_interconnect_1_position_y_s1_readdata),                  //                                                 .readdata
		.position_z_s1_address                                  (mm_interconnect_1_position_z_s1_address),                   //                                    position_z_s1.address
		.position_z_s1_readdata                                 (mm_interconnect_1_position_z_s1_readdata),                  //                                                 .readdata
		.settings_acceleration_e0_s1_address                    (mm_interconnect_1_settings_acceleration_e0_s1_address),     //                      settings_acceleration_e0_s1.address
		.settings_acceleration_e0_s1_write                      (mm_interconnect_1_settings_acceleration_e0_s1_write),       //                                                 .write
		.settings_acceleration_e0_s1_readdata                   (mm_interconnect_1_settings_acceleration_e0_s1_readdata),    //                                                 .readdata
		.settings_acceleration_e0_s1_writedata                  (mm_interconnect_1_settings_acceleration_e0_s1_writedata),   //                                                 .writedata
		.settings_acceleration_e0_s1_chipselect                 (mm_interconnect_1_settings_acceleration_e0_s1_chipselect),  //                                                 .chipselect
		.settings_acceleration_e1_s1_address                    (mm_interconnect_1_settings_acceleration_e1_s1_address),     //                      settings_acceleration_e1_s1.address
		.settings_acceleration_e1_s1_write                      (mm_interconnect_1_settings_acceleration_e1_s1_write),       //                                                 .write
		.settings_acceleration_e1_s1_readdata                   (mm_interconnect_1_settings_acceleration_e1_s1_readdata),    //                                                 .readdata
		.settings_acceleration_e1_s1_writedata                  (mm_interconnect_1_settings_acceleration_e1_s1_writedata),   //                                                 .writedata
		.settings_acceleration_e1_s1_chipselect                 (mm_interconnect_1_settings_acceleration_e1_s1_chipselect),  //                                                 .chipselect
		.settings_acceleration_x_s1_address                     (mm_interconnect_1_settings_acceleration_x_s1_address),      //                       settings_acceleration_x_s1.address
		.settings_acceleration_x_s1_write                       (mm_interconnect_1_settings_acceleration_x_s1_write),        //                                                 .write
		.settings_acceleration_x_s1_readdata                    (mm_interconnect_1_settings_acceleration_x_s1_readdata),     //                                                 .readdata
		.settings_acceleration_x_s1_writedata                   (mm_interconnect_1_settings_acceleration_x_s1_writedata),    //                                                 .writedata
		.settings_acceleration_x_s1_chipselect                  (mm_interconnect_1_settings_acceleration_x_s1_chipselect),   //                                                 .chipselect
		.settings_acceleration_y_s1_address                     (mm_interconnect_1_settings_acceleration_y_s1_address),      //                       settings_acceleration_y_s1.address
		.settings_acceleration_y_s1_write                       (mm_interconnect_1_settings_acceleration_y_s1_write),        //                                                 .write
		.settings_acceleration_y_s1_readdata                    (mm_interconnect_1_settings_acceleration_y_s1_readdata),     //                                                 .readdata
		.settings_acceleration_y_s1_writedata                   (mm_interconnect_1_settings_acceleration_y_s1_writedata),    //                                                 .writedata
		.settings_acceleration_y_s1_chipselect                  (mm_interconnect_1_settings_acceleration_y_s1_chipselect),   //                                                 .chipselect
		.settings_acceleration_z_s1_address                     (mm_interconnect_1_settings_acceleration_z_s1_address),      //                       settings_acceleration_z_s1.address
		.settings_acceleration_z_s1_write                       (mm_interconnect_1_settings_acceleration_z_s1_write),        //                                                 .write
		.settings_acceleration_z_s1_readdata                    (mm_interconnect_1_settings_acceleration_z_s1_readdata),     //                                                 .readdata
		.settings_acceleration_z_s1_writedata                   (mm_interconnect_1_settings_acceleration_z_s1_writedata),    //                                                 .writedata
		.settings_acceleration_z_s1_chipselect                  (mm_interconnect_1_settings_acceleration_z_s1_chipselect),   //                                                 .chipselect
		.settings_jerk_e0_s1_address                            (mm_interconnect_1_settings_jerk_e0_s1_address),             //                              settings_jerk_e0_s1.address
		.settings_jerk_e0_s1_write                              (mm_interconnect_1_settings_jerk_e0_s1_write),               //                                                 .write
		.settings_jerk_e0_s1_readdata                           (mm_interconnect_1_settings_jerk_e0_s1_readdata),            //                                                 .readdata
		.settings_jerk_e0_s1_writedata                          (mm_interconnect_1_settings_jerk_e0_s1_writedata),           //                                                 .writedata
		.settings_jerk_e0_s1_chipselect                         (mm_interconnect_1_settings_jerk_e0_s1_chipselect),          //                                                 .chipselect
		.settings_jerk_e1_s1_address                            (mm_interconnect_1_settings_jerk_e1_s1_address),             //                              settings_jerk_e1_s1.address
		.settings_jerk_e1_s1_write                              (mm_interconnect_1_settings_jerk_e1_s1_write),               //                                                 .write
		.settings_jerk_e1_s1_readdata                           (mm_interconnect_1_settings_jerk_e1_s1_readdata),            //                                                 .readdata
		.settings_jerk_e1_s1_writedata                          (mm_interconnect_1_settings_jerk_e1_s1_writedata),           //                                                 .writedata
		.settings_jerk_e1_s1_chipselect                         (mm_interconnect_1_settings_jerk_e1_s1_chipselect),          //                                                 .chipselect
		.settings_jerk_x_s1_address                             (mm_interconnect_1_settings_jerk_x_s1_address),              //                               settings_jerk_x_s1.address
		.settings_jerk_x_s1_write                               (mm_interconnect_1_settings_jerk_x_s1_write),                //                                                 .write
		.settings_jerk_x_s1_readdata                            (mm_interconnect_1_settings_jerk_x_s1_readdata),             //                                                 .readdata
		.settings_jerk_x_s1_writedata                           (mm_interconnect_1_settings_jerk_x_s1_writedata),            //                                                 .writedata
		.settings_jerk_x_s1_chipselect                          (mm_interconnect_1_settings_jerk_x_s1_chipselect),           //                                                 .chipselect
		.settings_jerk_y_s1_address                             (mm_interconnect_1_settings_jerk_y_s1_address),              //                               settings_jerk_y_s1.address
		.settings_jerk_y_s1_write                               (mm_interconnect_1_settings_jerk_y_s1_write),                //                                                 .write
		.settings_jerk_y_s1_readdata                            (mm_interconnect_1_settings_jerk_y_s1_readdata),             //                                                 .readdata
		.settings_jerk_y_s1_writedata                           (mm_interconnect_1_settings_jerk_y_s1_writedata),            //                                                 .writedata
		.settings_jerk_y_s1_chipselect                          (mm_interconnect_1_settings_jerk_y_s1_chipselect),           //                                                 .chipselect
		.settings_jerk_z_s1_address                             (mm_interconnect_1_settings_jerk_z_s1_address),              //                               settings_jerk_z_s1.address
		.settings_jerk_z_s1_write                               (mm_interconnect_1_settings_jerk_z_s1_write),                //                                                 .write
		.settings_jerk_z_s1_readdata                            (mm_interconnect_1_settings_jerk_z_s1_readdata),             //                                                 .readdata
		.settings_jerk_z_s1_writedata                           (mm_interconnect_1_settings_jerk_z_s1_writedata),            //                                                 .writedata
		.settings_jerk_z_s1_chipselect                          (mm_interconnect_1_settings_jerk_z_s1_chipselect),           //                                                 .chipselect
		.settings_max_speed_e0_s1_address                       (mm_interconnect_1_settings_max_speed_e0_s1_address),        //                         settings_max_speed_e0_s1.address
		.settings_max_speed_e0_s1_write                         (mm_interconnect_1_settings_max_speed_e0_s1_write),          //                                                 .write
		.settings_max_speed_e0_s1_readdata                      (mm_interconnect_1_settings_max_speed_e0_s1_readdata),       //                                                 .readdata
		.settings_max_speed_e0_s1_writedata                     (mm_interconnect_1_settings_max_speed_e0_s1_writedata),      //                                                 .writedata
		.settings_max_speed_e0_s1_chipselect                    (mm_interconnect_1_settings_max_speed_e0_s1_chipselect),     //                                                 .chipselect
		.settings_max_speed_e1_s1_address                       (mm_interconnect_1_settings_max_speed_e1_s1_address),        //                         settings_max_speed_e1_s1.address
		.settings_max_speed_e1_s1_write                         (mm_interconnect_1_settings_max_speed_e1_s1_write),          //                                                 .write
		.settings_max_speed_e1_s1_readdata                      (mm_interconnect_1_settings_max_speed_e1_s1_readdata),       //                                                 .readdata
		.settings_max_speed_e1_s1_writedata                     (mm_interconnect_1_settings_max_speed_e1_s1_writedata),      //                                                 .writedata
		.settings_max_speed_e1_s1_chipselect                    (mm_interconnect_1_settings_max_speed_e1_s1_chipselect),     //                                                 .chipselect
		.settings_max_speed_x_s1_address                        (mm_interconnect_1_settings_max_speed_x_s1_address),         //                          settings_max_speed_x_s1.address
		.settings_max_speed_x_s1_write                          (mm_interconnect_1_settings_max_speed_x_s1_write),           //                                                 .write
		.settings_max_speed_x_s1_readdata                       (mm_interconnect_1_settings_max_speed_x_s1_readdata),        //                                                 .readdata
		.settings_max_speed_x_s1_writedata                      (mm_interconnect_1_settings_max_speed_x_s1_writedata),       //                                                 .writedata
		.settings_max_speed_x_s1_chipselect                     (mm_interconnect_1_settings_max_speed_x_s1_chipselect),      //                                                 .chipselect
		.settings_max_speed_y_s1_address                        (mm_interconnect_1_settings_max_speed_y_s1_address),         //                          settings_max_speed_y_s1.address
		.settings_max_speed_y_s1_write                          (mm_interconnect_1_settings_max_speed_y_s1_write),           //                                                 .write
		.settings_max_speed_y_s1_readdata                       (mm_interconnect_1_settings_max_speed_y_s1_readdata),        //                                                 .readdata
		.settings_max_speed_y_s1_writedata                      (mm_interconnect_1_settings_max_speed_y_s1_writedata),       //                                                 .writedata
		.settings_max_speed_y_s1_chipselect                     (mm_interconnect_1_settings_max_speed_y_s1_chipselect),      //                                                 .chipselect
		.settings_max_speed_z_s1_address                        (mm_interconnect_1_settings_max_speed_z_s1_address),         //                          settings_max_speed_z_s1.address
		.settings_max_speed_z_s1_write                          (mm_interconnect_1_settings_max_speed_z_s1_write),           //                                                 .write
		.settings_max_speed_z_s1_readdata                       (mm_interconnect_1_settings_max_speed_z_s1_readdata),        //                                                 .readdata
		.settings_max_speed_z_s1_writedata                      (mm_interconnect_1_settings_max_speed_z_s1_writedata),       //                                                 .writedata
		.settings_max_speed_z_s1_chipselect                     (mm_interconnect_1_settings_max_speed_z_s1_chipselect),      //                                                 .chipselect
		.settings_max_temp_bed_s1_address                       (mm_interconnect_1_settings_max_temp_bed_s1_address),        //                         settings_max_temp_bed_s1.address
		.settings_max_temp_bed_s1_write                         (mm_interconnect_1_settings_max_temp_bed_s1_write),          //                                                 .write
		.settings_max_temp_bed_s1_readdata                      (mm_interconnect_1_settings_max_temp_bed_s1_readdata),       //                                                 .readdata
		.settings_max_temp_bed_s1_writedata                     (mm_interconnect_1_settings_max_temp_bed_s1_writedata),      //                                                 .writedata
		.settings_max_temp_bed_s1_chipselect                    (mm_interconnect_1_settings_max_temp_bed_s1_chipselect),     //                                                 .chipselect
		.settings_max_temp_e0_s1_address                        (mm_interconnect_1_settings_max_temp_e0_s1_address),         //                          settings_max_temp_e0_s1.address
		.settings_max_temp_e0_s1_write                          (mm_interconnect_1_settings_max_temp_e0_s1_write),           //                                                 .write
		.settings_max_temp_e0_s1_readdata                       (mm_interconnect_1_settings_max_temp_e0_s1_readdata),        //                                                 .readdata
		.settings_max_temp_e0_s1_writedata                      (mm_interconnect_1_settings_max_temp_e0_s1_writedata),       //                                                 .writedata
		.settings_max_temp_e0_s1_chipselect                     (mm_interconnect_1_settings_max_temp_e0_s1_chipselect),      //                                                 .chipselect
		.settings_max_temp_e1_s1_address                        (mm_interconnect_1_settings_max_temp_e1_s1_address),         //                          settings_max_temp_e1_s1.address
		.settings_max_temp_e1_s1_write                          (mm_interconnect_1_settings_max_temp_e1_s1_write),           //                                                 .write
		.settings_max_temp_e1_s1_readdata                       (mm_interconnect_1_settings_max_temp_e1_s1_readdata),        //                                                 .readdata
		.settings_max_temp_e1_s1_writedata                      (mm_interconnect_1_settings_max_temp_e1_s1_writedata),       //                                                 .writedata
		.settings_max_temp_e1_s1_chipselect                     (mm_interconnect_1_settings_max_temp_e1_s1_chipselect),      //                                                 .chipselect
		.step_e0_now_s1_address                                 (mm_interconnect_1_step_e0_now_s1_address),                  //                                   step_e0_now_s1.address
		.step_e0_now_s1_readdata                                (mm_interconnect_1_step_e0_now_s1_readdata),                 //                                                 .readdata
		.step_e1_now_s1_address                                 (mm_interconnect_1_step_e1_now_s1_address),                  //                                   step_e1_now_s1.address
		.step_e1_now_s1_readdata                                (mm_interconnect_1_step_e1_now_s1_readdata),                 //                                                 .readdata
		.step_x_now_s1_address                                  (mm_interconnect_1_step_x_now_s1_address),                   //                                    step_x_now_s1.address
		.step_x_now_s1_readdata                                 (mm_interconnect_1_step_x_now_s1_readdata),                  //                                                 .readdata
		.step_y_now_s1_address                                  (mm_interconnect_1_step_y_now_s1_address),                   //                                    step_y_now_s1.address
		.step_y_now_s1_readdata                                 (mm_interconnect_1_step_y_now_s1_readdata),                  //                                                 .readdata
		.step_z_now_s1_address                                  (mm_interconnect_1_step_z_now_s1_address),                   //                                    step_z_now_s1.address
		.step_z_now_s1_readdata                                 (mm_interconnect_1_step_z_now_s1_readdata),                  //                                                 .readdata
		.sysid_qsys_control_slave_address                       (mm_interconnect_1_sysid_qsys_control_slave_address),        //                         sysid_qsys_control_slave.address
		.sysid_qsys_control_slave_readdata                      (mm_interconnect_1_sysid_qsys_control_slave_readdata),       //                                                 .readdata
		.temp_0_s1_address                                      (mm_interconnect_1_temp_0_s1_address),                       //                                        temp_0_s1.address
		.temp_0_s1_readdata                                     (mm_interconnect_1_temp_0_s1_readdata),                      //                                                 .readdata
		.temp_1_s1_address                                      (mm_interconnect_1_temp_1_s1_address),                       //                                        temp_1_s1.address
		.temp_1_s1_readdata                                     (mm_interconnect_1_temp_1_s1_readdata),                      //                                                 .readdata
		.temp_2_s1_address                                      (mm_interconnect_1_temp_2_s1_address),                       //                                        temp_2_s1.address
		.temp_2_s1_readdata                                     (mm_interconnect_1_temp_2_s1_readdata),                      //                                                 .readdata
		.timing_e0_0_s1_address                                 (mm_interconnect_1_timing_e0_0_s1_address),                  //                                   timing_e0_0_s1.address
		.timing_e0_0_s1_readdata                                (mm_interconnect_1_timing_e0_0_s1_readdata),                 //                                                 .readdata
		.timing_e0_1_s1_address                                 (mm_interconnect_1_timing_e0_1_s1_address),                  //                                   timing_e0_1_s1.address
		.timing_e0_1_s1_readdata                                (mm_interconnect_1_timing_e0_1_s1_readdata),                 //                                                 .readdata
		.timing_e0_2_s1_address                                 (mm_interconnect_1_timing_e0_2_s1_address),                  //                                   timing_e0_2_s1.address
		.timing_e0_2_s1_readdata                                (mm_interconnect_1_timing_e0_2_s1_readdata),                 //                                                 .readdata
		.timing_e0_3_s1_address                                 (mm_interconnect_1_timing_e0_3_s1_address),                  //                                   timing_e0_3_s1.address
		.timing_e0_3_s1_readdata                                (mm_interconnect_1_timing_e0_3_s1_readdata),                 //                                                 .readdata
		.timing_e1_0_s1_address                                 (mm_interconnect_1_timing_e1_0_s1_address),                  //                                   timing_e1_0_s1.address
		.timing_e1_0_s1_readdata                                (mm_interconnect_1_timing_e1_0_s1_readdata),                 //                                                 .readdata
		.timing_e1_1_s1_address                                 (mm_interconnect_1_timing_e1_1_s1_address),                  //                                   timing_e1_1_s1.address
		.timing_e1_1_s1_readdata                                (mm_interconnect_1_timing_e1_1_s1_readdata),                 //                                                 .readdata
		.timing_e1_2_s1_address                                 (mm_interconnect_1_timing_e1_2_s1_address),                  //                                   timing_e1_2_s1.address
		.timing_e1_2_s1_readdata                                (mm_interconnect_1_timing_e1_2_s1_readdata),                 //                                                 .readdata
		.timing_e1_3_s1_address                                 (mm_interconnect_1_timing_e1_3_s1_address),                  //                                   timing_e1_3_s1.address
		.timing_e1_3_s1_readdata                                (mm_interconnect_1_timing_e1_3_s1_readdata),                 //                                                 .readdata
		.timing_x_0_s1_address                                  (mm_interconnect_1_timing_x_0_s1_address),                   //                                    timing_x_0_s1.address
		.timing_x_0_s1_readdata                                 (mm_interconnect_1_timing_x_0_s1_readdata),                  //                                                 .readdata
		.timing_x_1_s1_address                                  (mm_interconnect_1_timing_x_1_s1_address),                   //                                    timing_x_1_s1.address
		.timing_x_1_s1_readdata                                 (mm_interconnect_1_timing_x_1_s1_readdata),                  //                                                 .readdata
		.timing_x_2_s1_address                                  (mm_interconnect_1_timing_x_2_s1_address),                   //                                    timing_x_2_s1.address
		.timing_x_2_s1_readdata                                 (mm_interconnect_1_timing_x_2_s1_readdata),                  //                                                 .readdata
		.timing_x_3_s1_address                                  (mm_interconnect_1_timing_x_3_s1_address),                   //                                    timing_x_3_s1.address
		.timing_x_3_s1_readdata                                 (mm_interconnect_1_timing_x_3_s1_readdata),                  //                                                 .readdata
		.timing_y_0_s1_address                                  (mm_interconnect_1_timing_y_0_s1_address),                   //                                    timing_y_0_s1.address
		.timing_y_0_s1_readdata                                 (mm_interconnect_1_timing_y_0_s1_readdata),                  //                                                 .readdata
		.timing_y_1_s1_address                                  (mm_interconnect_1_timing_y_1_s1_address),                   //                                    timing_y_1_s1.address
		.timing_y_1_s1_readdata                                 (mm_interconnect_1_timing_y_1_s1_readdata),                  //                                                 .readdata
		.timing_y_2_s1_address                                  (mm_interconnect_1_timing_y_2_s1_address),                   //                                    timing_y_2_s1.address
		.timing_y_2_s1_readdata                                 (mm_interconnect_1_timing_y_2_s1_readdata),                  //                                                 .readdata
		.timing_y_3_s1_address                                  (mm_interconnect_1_timing_y_3_s1_address),                   //                                    timing_y_3_s1.address
		.timing_y_3_s1_readdata                                 (mm_interconnect_1_timing_y_3_s1_readdata),                  //                                                 .readdata
		.timing_z_0_s1_address                                  (mm_interconnect_1_timing_z_0_s1_address),                   //                                    timing_z_0_s1.address
		.timing_z_0_s1_readdata                                 (mm_interconnect_1_timing_z_0_s1_readdata),                  //                                                 .readdata
		.timing_z_1_s1_address                                  (mm_interconnect_1_timing_z_1_s1_address),                   //                                    timing_z_1_s1.address
		.timing_z_1_s1_readdata                                 (mm_interconnect_1_timing_z_1_s1_readdata),                  //                                                 .readdata
		.timing_z_2_s1_address                                  (mm_interconnect_1_timing_z_2_s1_address),                   //                                    timing_z_2_s1.address
		.timing_z_2_s1_readdata                                 (mm_interconnect_1_timing_z_2_s1_readdata),                  //                                                 .readdata
		.timing_z_3_s1_address                                  (mm_interconnect_1_timing_z_3_s1_address),                   //                                    timing_z_3_s1.address
		.timing_z_3_s1_readdata                                 (mm_interconnect_1_timing_z_3_s1_readdata)                   //                                                 .readdata
	);

	soc_system_mm_interconnect_2 mm_interconnect_2 (
		.hps_0_f2h_axi_slave_awid                                            (mm_interconnect_2_hps_0_f2h_axi_slave_awid),    //                                           hps_0_f2h_axi_slave.awid
		.hps_0_f2h_axi_slave_awaddr                                          (mm_interconnect_2_hps_0_f2h_axi_slave_awaddr),  //                                                              .awaddr
		.hps_0_f2h_axi_slave_awlen                                           (mm_interconnect_2_hps_0_f2h_axi_slave_awlen),   //                                                              .awlen
		.hps_0_f2h_axi_slave_awsize                                          (mm_interconnect_2_hps_0_f2h_axi_slave_awsize),  //                                                              .awsize
		.hps_0_f2h_axi_slave_awburst                                         (mm_interconnect_2_hps_0_f2h_axi_slave_awburst), //                                                              .awburst
		.hps_0_f2h_axi_slave_awlock                                          (mm_interconnect_2_hps_0_f2h_axi_slave_awlock),  //                                                              .awlock
		.hps_0_f2h_axi_slave_awcache                                         (mm_interconnect_2_hps_0_f2h_axi_slave_awcache), //                                                              .awcache
		.hps_0_f2h_axi_slave_awprot                                          (mm_interconnect_2_hps_0_f2h_axi_slave_awprot),  //                                                              .awprot
		.hps_0_f2h_axi_slave_awuser                                          (mm_interconnect_2_hps_0_f2h_axi_slave_awuser),  //                                                              .awuser
		.hps_0_f2h_axi_slave_awvalid                                         (mm_interconnect_2_hps_0_f2h_axi_slave_awvalid), //                                                              .awvalid
		.hps_0_f2h_axi_slave_awready                                         (mm_interconnect_2_hps_0_f2h_axi_slave_awready), //                                                              .awready
		.hps_0_f2h_axi_slave_wid                                             (mm_interconnect_2_hps_0_f2h_axi_slave_wid),     //                                                              .wid
		.hps_0_f2h_axi_slave_wdata                                           (mm_interconnect_2_hps_0_f2h_axi_slave_wdata),   //                                                              .wdata
		.hps_0_f2h_axi_slave_wstrb                                           (mm_interconnect_2_hps_0_f2h_axi_slave_wstrb),   //                                                              .wstrb
		.hps_0_f2h_axi_slave_wlast                                           (mm_interconnect_2_hps_0_f2h_axi_slave_wlast),   //                                                              .wlast
		.hps_0_f2h_axi_slave_wvalid                                          (mm_interconnect_2_hps_0_f2h_axi_slave_wvalid),  //                                                              .wvalid
		.hps_0_f2h_axi_slave_wready                                          (mm_interconnect_2_hps_0_f2h_axi_slave_wready),  //                                                              .wready
		.hps_0_f2h_axi_slave_bid                                             (mm_interconnect_2_hps_0_f2h_axi_slave_bid),     //                                                              .bid
		.hps_0_f2h_axi_slave_bresp                                           (mm_interconnect_2_hps_0_f2h_axi_slave_bresp),   //                                                              .bresp
		.hps_0_f2h_axi_slave_bvalid                                          (mm_interconnect_2_hps_0_f2h_axi_slave_bvalid),  //                                                              .bvalid
		.hps_0_f2h_axi_slave_bready                                          (mm_interconnect_2_hps_0_f2h_axi_slave_bready),  //                                                              .bready
		.hps_0_f2h_axi_slave_arid                                            (mm_interconnect_2_hps_0_f2h_axi_slave_arid),    //                                                              .arid
		.hps_0_f2h_axi_slave_araddr                                          (mm_interconnect_2_hps_0_f2h_axi_slave_araddr),  //                                                              .araddr
		.hps_0_f2h_axi_slave_arlen                                           (mm_interconnect_2_hps_0_f2h_axi_slave_arlen),   //                                                              .arlen
		.hps_0_f2h_axi_slave_arsize                                          (mm_interconnect_2_hps_0_f2h_axi_slave_arsize),  //                                                              .arsize
		.hps_0_f2h_axi_slave_arburst                                         (mm_interconnect_2_hps_0_f2h_axi_slave_arburst), //                                                              .arburst
		.hps_0_f2h_axi_slave_arlock                                          (mm_interconnect_2_hps_0_f2h_axi_slave_arlock),  //                                                              .arlock
		.hps_0_f2h_axi_slave_arcache                                         (mm_interconnect_2_hps_0_f2h_axi_slave_arcache), //                                                              .arcache
		.hps_0_f2h_axi_slave_arprot                                          (mm_interconnect_2_hps_0_f2h_axi_slave_arprot),  //                                                              .arprot
		.hps_0_f2h_axi_slave_aruser                                          (mm_interconnect_2_hps_0_f2h_axi_slave_aruser),  //                                                              .aruser
		.hps_0_f2h_axi_slave_arvalid                                         (mm_interconnect_2_hps_0_f2h_axi_slave_arvalid), //                                                              .arvalid
		.hps_0_f2h_axi_slave_arready                                         (mm_interconnect_2_hps_0_f2h_axi_slave_arready), //                                                              .arready
		.hps_0_f2h_axi_slave_rid                                             (mm_interconnect_2_hps_0_f2h_axi_slave_rid),     //                                                              .rid
		.hps_0_f2h_axi_slave_rdata                                           (mm_interconnect_2_hps_0_f2h_axi_slave_rdata),   //                                                              .rdata
		.hps_0_f2h_axi_slave_rresp                                           (mm_interconnect_2_hps_0_f2h_axi_slave_rresp),   //                                                              .rresp
		.hps_0_f2h_axi_slave_rlast                                           (mm_interconnect_2_hps_0_f2h_axi_slave_rlast),   //                                                              .rlast
		.hps_0_f2h_axi_slave_rvalid                                          (mm_interconnect_2_hps_0_f2h_axi_slave_rvalid),  //                                                              .rvalid
		.hps_0_f2h_axi_slave_rready                                          (mm_interconnect_2_hps_0_f2h_axi_slave_rready),  //                                                              .rready
		.clk_0_clk_clk                                                       (clk_clk),                                       //                                                     clk_0_clk.clk
		.hps_0_f2h_axi_slave_agent_reset_sink_reset_bridge_in_reset_reset    (rst_controller_001_reset_out_reset),            //    hps_0_f2h_axi_slave_agent_reset_sink_reset_bridge_in_reset.reset
		.hps_only_master_clk_reset_reset_bridge_in_reset_reset               (rst_controller_reset_out_reset),                //               hps_only_master_clk_reset_reset_bridge_in_reset.reset
		.hps_only_master_master_translator_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                // hps_only_master_master_translator_reset_reset_bridge_in_reset.reset
		.hps_only_master_master_address                                      (hps_only_master_master_address),                //                                        hps_only_master_master.address
		.hps_only_master_master_waitrequest                                  (hps_only_master_master_waitrequest),            //                                                              .waitrequest
		.hps_only_master_master_byteenable                                   (hps_only_master_master_byteenable),             //                                                              .byteenable
		.hps_only_master_master_read                                         (hps_only_master_master_read),                   //                                                              .read
		.hps_only_master_master_readdata                                     (hps_only_master_master_readdata),               //                                                              .readdata
		.hps_only_master_master_readdatavalid                                (hps_only_master_master_readdatavalid),          //                                                              .readdatavalid
		.hps_only_master_master_write                                        (hps_only_master_master_write),                  //                                                              .write
		.hps_only_master_master_writedata                                    (hps_only_master_master_writedata)               //                                                              .writedata
	);

	soc_system_mm_interconnect_3 mm_interconnect_3 (
		.clk_0_clk_clk                                                           (clk_clk),                                               //                                                         clk_0_clk.clk
		.f2sdram_only_master_clk_reset_reset_bridge_in_reset_reset               (rst_controller_reset_out_reset),                        //               f2sdram_only_master_clk_reset_reset_bridge_in_reset.reset
		.f2sdram_only_master_master_translator_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                        // f2sdram_only_master_master_translator_reset_reset_bridge_in_reset.reset
		.hps_0_f2h_sdram0_data_translator_reset_reset_bridge_in_reset_reset      (rst_controller_001_reset_out_reset),                    //      hps_0_f2h_sdram0_data_translator_reset_reset_bridge_in_reset.reset
		.f2sdram_only_master_master_address                                      (f2sdram_only_master_master_address),                    //                                        f2sdram_only_master_master.address
		.f2sdram_only_master_master_waitrequest                                  (f2sdram_only_master_master_waitrequest),                //                                                                  .waitrequest
		.f2sdram_only_master_master_byteenable                                   (f2sdram_only_master_master_byteenable),                 //                                                                  .byteenable
		.f2sdram_only_master_master_read                                         (f2sdram_only_master_master_read),                       //                                                                  .read
		.f2sdram_only_master_master_readdata                                     (f2sdram_only_master_master_readdata),                   //                                                                  .readdata
		.f2sdram_only_master_master_readdatavalid                                (f2sdram_only_master_master_readdatavalid),              //                                                                  .readdatavalid
		.f2sdram_only_master_master_write                                        (f2sdram_only_master_master_write),                      //                                                                  .write
		.f2sdram_only_master_master_writedata                                    (f2sdram_only_master_master_writedata),                  //                                                                  .writedata
		.hps_0_f2h_sdram0_data_address                                           (mm_interconnect_3_hps_0_f2h_sdram0_data_address),       //                                             hps_0_f2h_sdram0_data.address
		.hps_0_f2h_sdram0_data_write                                             (mm_interconnect_3_hps_0_f2h_sdram0_data_write),         //                                                                  .write
		.hps_0_f2h_sdram0_data_read                                              (mm_interconnect_3_hps_0_f2h_sdram0_data_read),          //                                                                  .read
		.hps_0_f2h_sdram0_data_readdata                                          (mm_interconnect_3_hps_0_f2h_sdram0_data_readdata),      //                                                                  .readdata
		.hps_0_f2h_sdram0_data_writedata                                         (mm_interconnect_3_hps_0_f2h_sdram0_data_writedata),     //                                                                  .writedata
		.hps_0_f2h_sdram0_data_burstcount                                        (mm_interconnect_3_hps_0_f2h_sdram0_data_burstcount),    //                                                                  .burstcount
		.hps_0_f2h_sdram0_data_byteenable                                        (mm_interconnect_3_hps_0_f2h_sdram0_data_byteenable),    //                                                                  .byteenable
		.hps_0_f2h_sdram0_data_readdatavalid                                     (mm_interconnect_3_hps_0_f2h_sdram0_data_readdatavalid), //                                                                  .readdatavalid
		.hps_0_f2h_sdram0_data_waitrequest                                       (mm_interconnect_3_hps_0_f2h_sdram0_data_waitrequest)    //                                                                  .waitrequest
	);

	soc_system_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (ilc_irq_irq)                     //    sender.irq
	);

	soc_system_irq_mapper_001 irq_mapper_001 (
		.clk           (),                         //       clk.clk
		.reset         (),                         // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq), // receiver0.irq
		.sender_irq    (hps_0_f2h_irq0_irq)        //    sender.irq
	);

	soc_system_irq_mapper_002 irq_mapper_002 (
		.clk        (),                   //       clk.clk
		.reset      (),                   // clk_reset.reset
		.sender_irq (hps_0_f2h_irq1_irq)  //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~hps_0_h2f_reset_reset_n),           // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
